//systemVerilog HDL for "MAD_RISC_tb", "REGFILE_tb" "systemVerilog"


module REGFILE_tb ( );

endmodule
