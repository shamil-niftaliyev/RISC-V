 module SINGLECORE (
	CLK, 
	RST, 
	INSTR, 
	DMEMRD, 
	PC, 
	ALURSLT, 
	WRDATA, 
	MEMWRITE);
   input CLK;
   input RST;
   input [31:0] INSTR;
   input [31:0] DMEMRD;
   output [31:0] PC;
   output [31:0] ALURSLT;
   output [31:0] WRDATA;
   output MEMWRITE;

   // Internal wires
   wire FE_PDN1444_FE_OFN34_n_1383;
   wire FE_PDN1443_FE_OFN34_n_1383;
   wire FE_OFN1442_n_111;
   wire FE_OFN1441_n_2619;
   wire CTS_61;
   wire CTS_60;
   wire CTS_7;
   wire CTS_6;
   wire CTS_5;
   wire CTS_4;
   wire CTS_3;
   wire CTS_2;
   wire CTS_1;
   wire CTS_9;
   wire CTS_59;
   wire CTS_58;
   wire CTS_57;
   wire CTS_56;
   wire CTS_55;
   wire CTS_54;
   wire CTS_53;
   wire CTS_52;
   wire CTS_51;
   wire CTS_25;
   wire CTS_24;
   wire CTS_23;
   wire CTS_27;
   wire CTS_50;
   wire CTS_49;
   wire CTS_48;
   wire CTS_47;
   wire CTS_46;
   wire CTS_45;
   wire CTS_44;
   wire CTS_43;
   wire CTS_42;
   wire CTS_20;
   wire CTS_19;
   wire CTS_18;
   wire CTS_17;
   wire CTS_16;
   wire CTS_15;
   wire CTS_22;
   wire CTS_41;
   wire CTS_12;
   wire CTS_11;
   wire CTS_10;
   wire CTS_14;
   wire CTS_40;
   wire CTS_39;
   wire CTS_38;
   wire CTS_37;
   wire CTS_36;
   wire CTS_35;
   wire CTS_34;
   wire CTS_33;
   wire CTS_32;
   wire CTS_31;
   wire CTS_30;
   wire CTS_29;
   wire CTS_28;
   wire CTS_26;
   wire CTS_21;
   wire CTS_13;
   wire CTS_8;
   wire FE_OFN119_n_95;
   wire FE_OFN118_n_1198;
   wire FE_OFN117_n_154;
   wire FE_OFN116_n_152;
   wire FE_OFN115_n_152;
   wire FE_OFN114_n_150;
   wire FE_OFN113_n_148;
   wire FE_OFN112_n_146;
   wire FE_OFN111_n_144;
   wire FE_OFN110_n_142;
   wire FE_OFN109_n_142;
   wire FE_OFN108_n_140;
   wire FE_OFN107_n_138;
   wire FE_OFN106_n_136;
   wire FE_OFN105_n_134;
   wire FE_OFN104_n_134;
   wire FE_OFN103_n_132;
   wire FE_OFN102_n_130;
   wire FE_OFN101_n_128;
   wire FE_OFN100_n_127;
   wire FE_OFN99_n_125;
   wire FE_OFN98_n_125;
   wire FE_OFN97_n_123;
   wire FE_OFN96_n_121;
   wire FE_OFN95_n_119;
   wire FE_OFN94_n_119;
   wire FE_OFN93_n_117;
   wire FE_OFN92_n_115;
   wire FE_OFN91_n_113;
   wire FE_OFN90_n_111;
   wire FE_OFN89_n_109;
   wire FE_OFN88_n_107;
   wire FE_OFN87_n_105;
   wire FE_OFN86_n_103;
   wire FE_OFN85_n_101;
   wire FE_OFN84_n_99;
   wire FE_OFN83_n_97;
   wire FE_OFN82_n_93;
   wire FE_OFN81_n_86;
   wire FE_OFN80_n_85;
   wire FE_OFN79_n_82;
   wire FE_OFN78_n_79;
   wire FE_OFN77_n_76;
   wire FE_OFN76_n_75;
   wire FE_OFN75_n_73;
   wire FE_OFN74_n_72;
   wire FE_OFN73_n_1449;
   wire FE_OFN72_n_1448;
   wire FE_OFN69_n_1443;
   wire FE_OFN68_n_1442;
   wire FE_OFN67_n_1441;
   wire FE_OFN66_n_1440;
   wire FE_OFN65_n_1438;
   wire FE_OFN64_n_1436;
   wire FE_OFN63_n_1432;
   wire FE_OFN62_n_1429;
   wire FE_OFN60_n_1425;
   wire FE_OFN59_n_1423;
   wire FE_OFN58_n_1422;
   wire FE_OFN57_n_1419;
   wire FE_OFN56_n_1415;
   wire FE_OFN55_n_1413;
   wire FE_OFN54_n_1411;
   wire FE_OFN53_n_1409;
   wire FE_OFN52_n_1408;
   wire FE_OFN49_n_1404;
   wire FE_OFN48_n_1401;
   wire FE_OFN47_n_1400;
   wire FE_OFN46_n_1398;
   wire FE_OFN45_n_1397;
   wire FE_OFN44_n_1396;
   wire FE_OFN43_n_1395;
   wire FE_OFN42_n_1393;
   wire FE_OFN41_n_1392;
   wire FE_OFN40_n_1391;
   wire FE_OFN39_n_1390;
   wire FE_OFN38_n_1389;
   wire FE_OFN36_n_1386;
   wire FE_OFN35_n_1385;
   wire FE_OFN34_n_1383;
   wire FE_OFN33_n_1381;
   wire FE_OFN32_n_1380;
   wire FE_OFN31_n_1379;
   wire FE_OFN29_n_1377;
   wire FE_OFN28_n_1376;
   wire FE_OFN27_n_1374;
   wire FE_OFN26_n_1371;
   wire FE_OFN25_n_1331;
   wire FE_OFN24_n_1162;
   wire FE_OFN23_n_91;
   wire FE_OFN22_n_90;
   wire FE_OFN21_n_89;
   wire FE_OFN19_n_88;
   wire FE_OFN17_n_87;
   wire FE_OFN16_n_84;
   wire FE_OFN15_n_83;
   wire FE_OFN13_n_80;
   wire FE_OFN12_n_78;
   wire FE_OFN10_n_77;
   wire FE_OFN9_n_74;
   wire FE_OFN8_n_71;
   wire FE_OFN6_n_70;
   wire FE_OFN5_n_69;
   wire FE_OFN4_n_67;
   wire FE_OFN3_n_64;
   wire FE_OFN2_n_62;
   wire FE_OFN0_n_2;
   wire DPATH_ADDBRANCH_add_422_17_n_596;
   wire DPATH_ADDBRANCH_add_422_17_n_599;
   wire DPATH_ADDBRANCH_add_422_17_n_601;
   wire DPATH_ADDBRANCH_add_422_17_n_603;
   wire DPATH_ADDBRANCH_add_422_17_n_605;
   wire DPATH_ADDBRANCH_add_422_17_n_607;
   wire DPATH_ADDBRANCH_add_422_17_n_609;
   wire DPATH_ADDBRANCH_add_422_17_n_611;
   wire DPATH_ADDBRANCH_add_422_17_n_613;
   wire DPATH_ADDBRANCH_add_422_17_n_615;
   wire DPATH_ADDBRANCH_add_422_17_n_617;
   wire DPATH_ADDBRANCH_add_422_17_n_619;
   wire DPATH_ADDBRANCH_add_422_17_n_621;
   wire DPATH_ADDBRANCH_add_422_17_n_623;
   wire DPATH_ADDBRANCH_add_422_17_n_625;
   wire DPATH_ADDBRANCH_add_422_17_n_627;
   wire DPATH_ADDBRANCH_add_422_17_n_629;
   wire DPATH_ADDBRANCH_add_422_17_n_631;
   wire DPATH_ADDBRANCH_add_422_17_n_633;
   wire DPATH_ADDBRANCH_add_422_17_n_635;
   wire DPATH_ADDBRANCH_add_422_17_n_637;
   wire DPATH_ADDBRANCH_add_422_17_n_639;
   wire DPATH_ADDBRANCH_add_422_17_n_641;
   wire DPATH_ADDBRANCH_add_422_17_n_643;
   wire DPATH_ADDBRANCH_add_422_17_n_645;
   wire DPATH_ADDBRANCH_add_422_17_n_647;
   wire DPATH_ADDBRANCH_add_422_17_n_649;
   wire DPATH_ADDBRANCH_add_422_17_n_651;
   wire DPATH_ADDBRANCH_add_422_17_n_653;
   wire DPATH_ADDBRANCH_add_422_17_n_655;
   wire DPATH_ADDFOUR_add_172_17_n_635;
   wire DPATH_ADDFOUR_add_172_17_n_637;
   wire DPATH_ADDFOUR_add_172_17_n_639;
   wire DPATH_ADDFOUR_add_172_17_n_641;
   wire DPATH_ADDFOUR_add_172_17_n_643;
   wire DPATH_ADDFOUR_add_172_17_n_645;
   wire DPATH_ADDFOUR_add_172_17_n_647;
   wire DPATH_ADDFOUR_add_172_17_n_649;
   wire DPATH_ADDFOUR_add_172_17_n_651;
   wire DPATH_ADDFOUR_add_172_17_n_653;
   wire DPATH_ADDFOUR_add_172_17_n_655;
   wire DPATH_ADDFOUR_add_172_17_n_657;
   wire DPATH_ADDFOUR_add_172_17_n_659;
   wire DPATH_ADDFOUR_add_172_17_n_661;
   wire DPATH_ADDFOUR_add_172_17_n_663;
   wire DPATH_ADDFOUR_add_172_17_n_665;
   wire DPATH_ADDFOUR_add_172_17_n_667;
   wire DPATH_ADDFOUR_add_172_17_n_669;
   wire DPATH_ADDFOUR_add_172_17_n_671;
   wire DPATH_ADDFOUR_add_172_17_n_673;
   wire DPATH_ADDFOUR_add_172_17_n_675;
   wire DPATH_ADDFOUR_add_172_17_n_677;
   wire DPATH_ADDFOUR_add_172_17_n_679;
   wire DPATH_ADDFOUR_add_172_17_n_681;
   wire DPATH_ADDFOUR_add_172_17_n_683;
   wire DPATH_ADDFOUR_add_172_17_n_685;
   wire DPATH_ADDFOUR_add_172_17_n_687;
   wire DPATH_ADDFOUR_add_172_17_n_689;
   wire DPATH_ALU_SUM_31__624;
   wire DPATH_A_31_;
   wire DPATH_B_31_;
   wire DPATH_RF_MEMORY_1__0_;
   wire DPATH_RF_MEMORY_1__1_;
   wire DPATH_RF_MEMORY_1__2_;
   wire DPATH_RF_MEMORY_1__3_;
   wire DPATH_RF_MEMORY_1__4_;
   wire DPATH_RF_MEMORY_1__5_;
   wire DPATH_RF_MEMORY_1__6_;
   wire DPATH_RF_MEMORY_1__7_;
   wire DPATH_RF_MEMORY_1__8_;
   wire DPATH_RF_MEMORY_1__9_;
   wire DPATH_RF_MEMORY_1__10_;
   wire DPATH_RF_MEMORY_1__11_;
   wire DPATH_RF_MEMORY_1__12_;
   wire DPATH_RF_MEMORY_1__13_;
   wire DPATH_RF_MEMORY_1__14_;
   wire DPATH_RF_MEMORY_1__15_;
   wire DPATH_RF_MEMORY_1__16_;
   wire DPATH_RF_MEMORY_1__17_;
   wire DPATH_RF_MEMORY_1__18_;
   wire DPATH_RF_MEMORY_1__19_;
   wire DPATH_RF_MEMORY_1__20_;
   wire DPATH_RF_MEMORY_1__21_;
   wire DPATH_RF_MEMORY_1__22_;
   wire DPATH_RF_MEMORY_1__23_;
   wire DPATH_RF_MEMORY_1__24_;
   wire DPATH_RF_MEMORY_1__25_;
   wire DPATH_RF_MEMORY_1__26_;
   wire DPATH_RF_MEMORY_1__27_;
   wire DPATH_RF_MEMORY_1__28_;
   wire DPATH_RF_MEMORY_1__29_;
   wire DPATH_RF_MEMORY_1__30_;
   wire DPATH_RF_MEMORY_1__31_;
   wire DPATH_RF_MEMORY_2__0_;
   wire DPATH_RF_MEMORY_2__1_;
   wire DPATH_RF_MEMORY_2__2_;
   wire DPATH_RF_MEMORY_2__3_;
   wire DPATH_RF_MEMORY_2__4_;
   wire DPATH_RF_MEMORY_2__5_;
   wire DPATH_RF_MEMORY_2__6_;
   wire DPATH_RF_MEMORY_2__7_;
   wire DPATH_RF_MEMORY_2__8_;
   wire DPATH_RF_MEMORY_2__9_;
   wire DPATH_RF_MEMORY_2__10_;
   wire DPATH_RF_MEMORY_2__11_;
   wire DPATH_RF_MEMORY_2__12_;
   wire DPATH_RF_MEMORY_2__13_;
   wire DPATH_RF_MEMORY_2__14_;
   wire DPATH_RF_MEMORY_2__15_;
   wire DPATH_RF_MEMORY_2__16_;
   wire DPATH_RF_MEMORY_2__17_;
   wire DPATH_RF_MEMORY_2__18_;
   wire DPATH_RF_MEMORY_2__19_;
   wire DPATH_RF_MEMORY_2__20_;
   wire DPATH_RF_MEMORY_2__21_;
   wire DPATH_RF_MEMORY_2__22_;
   wire DPATH_RF_MEMORY_2__23_;
   wire DPATH_RF_MEMORY_2__24_;
   wire DPATH_RF_MEMORY_2__25_;
   wire DPATH_RF_MEMORY_2__26_;
   wire DPATH_RF_MEMORY_2__27_;
   wire DPATH_RF_MEMORY_2__28_;
   wire DPATH_RF_MEMORY_2__29_;
   wire DPATH_RF_MEMORY_2__30_;
   wire DPATH_RF_MEMORY_2__31_;
   wire DPATH_RF_MEMORY_3__0_;
   wire DPATH_RF_MEMORY_3__1_;
   wire DPATH_RF_MEMORY_3__2_;
   wire DPATH_RF_MEMORY_3__3_;
   wire DPATH_RF_MEMORY_3__4_;
   wire DPATH_RF_MEMORY_3__5_;
   wire DPATH_RF_MEMORY_3__6_;
   wire DPATH_RF_MEMORY_3__7_;
   wire DPATH_RF_MEMORY_3__8_;
   wire DPATH_RF_MEMORY_3__9_;
   wire DPATH_RF_MEMORY_3__10_;
   wire DPATH_RF_MEMORY_3__11_;
   wire DPATH_RF_MEMORY_3__12_;
   wire DPATH_RF_MEMORY_3__13_;
   wire DPATH_RF_MEMORY_3__14_;
   wire DPATH_RF_MEMORY_3__15_;
   wire DPATH_RF_MEMORY_3__16_;
   wire DPATH_RF_MEMORY_3__17_;
   wire DPATH_RF_MEMORY_3__18_;
   wire DPATH_RF_MEMORY_3__19_;
   wire DPATH_RF_MEMORY_3__20_;
   wire DPATH_RF_MEMORY_3__21_;
   wire DPATH_RF_MEMORY_3__22_;
   wire DPATH_RF_MEMORY_3__23_;
   wire DPATH_RF_MEMORY_3__24_;
   wire DPATH_RF_MEMORY_3__25_;
   wire DPATH_RF_MEMORY_3__26_;
   wire DPATH_RF_MEMORY_3__27_;
   wire DPATH_RF_MEMORY_3__28_;
   wire DPATH_RF_MEMORY_3__29_;
   wire DPATH_RF_MEMORY_3__30_;
   wire DPATH_RF_MEMORY_3__31_;
   wire DPATH_RF_MEMORY_4__0_;
   wire DPATH_RF_MEMORY_4__1_;
   wire DPATH_RF_MEMORY_4__2_;
   wire DPATH_RF_MEMORY_4__3_;
   wire DPATH_RF_MEMORY_4__4_;
   wire DPATH_RF_MEMORY_4__5_;
   wire DPATH_RF_MEMORY_4__6_;
   wire DPATH_RF_MEMORY_4__7_;
   wire DPATH_RF_MEMORY_4__8_;
   wire DPATH_RF_MEMORY_4__9_;
   wire DPATH_RF_MEMORY_4__10_;
   wire DPATH_RF_MEMORY_4__11_;
   wire DPATH_RF_MEMORY_4__12_;
   wire DPATH_RF_MEMORY_4__13_;
   wire DPATH_RF_MEMORY_4__14_;
   wire DPATH_RF_MEMORY_4__15_;
   wire DPATH_RF_MEMORY_4__16_;
   wire DPATH_RF_MEMORY_4__17_;
   wire DPATH_RF_MEMORY_4__18_;
   wire DPATH_RF_MEMORY_4__19_;
   wire DPATH_RF_MEMORY_4__20_;
   wire DPATH_RF_MEMORY_4__21_;
   wire DPATH_RF_MEMORY_4__22_;
   wire DPATH_RF_MEMORY_4__23_;
   wire DPATH_RF_MEMORY_4__24_;
   wire DPATH_RF_MEMORY_4__25_;
   wire DPATH_RF_MEMORY_4__26_;
   wire DPATH_RF_MEMORY_4__27_;
   wire DPATH_RF_MEMORY_4__28_;
   wire DPATH_RF_MEMORY_4__29_;
   wire DPATH_RF_MEMORY_4__30_;
   wire DPATH_RF_MEMORY_4__31_;
   wire DPATH_RF_MEMORY_5__0_;
   wire DPATH_RF_MEMORY_5__1_;
   wire DPATH_RF_MEMORY_5__2_;
   wire DPATH_RF_MEMORY_5__3_;
   wire DPATH_RF_MEMORY_5__4_;
   wire DPATH_RF_MEMORY_5__5_;
   wire DPATH_RF_MEMORY_5__6_;
   wire DPATH_RF_MEMORY_5__7_;
   wire DPATH_RF_MEMORY_5__8_;
   wire DPATH_RF_MEMORY_5__9_;
   wire DPATH_RF_MEMORY_5__10_;
   wire DPATH_RF_MEMORY_5__11_;
   wire DPATH_RF_MEMORY_5__12_;
   wire DPATH_RF_MEMORY_5__13_;
   wire DPATH_RF_MEMORY_5__14_;
   wire DPATH_RF_MEMORY_5__15_;
   wire DPATH_RF_MEMORY_5__16_;
   wire DPATH_RF_MEMORY_5__17_;
   wire DPATH_RF_MEMORY_5__18_;
   wire DPATH_RF_MEMORY_5__19_;
   wire DPATH_RF_MEMORY_5__20_;
   wire DPATH_RF_MEMORY_5__21_;
   wire DPATH_RF_MEMORY_5__22_;
   wire DPATH_RF_MEMORY_5__23_;
   wire DPATH_RF_MEMORY_5__24_;
   wire DPATH_RF_MEMORY_5__25_;
   wire DPATH_RF_MEMORY_5__26_;
   wire DPATH_RF_MEMORY_5__27_;
   wire DPATH_RF_MEMORY_5__28_;
   wire DPATH_RF_MEMORY_5__29_;
   wire DPATH_RF_MEMORY_5__30_;
   wire DPATH_RF_MEMORY_5__31_;
   wire DPATH_RF_MEMORY_6__0_;
   wire DPATH_RF_MEMORY_6__1_;
   wire DPATH_RF_MEMORY_6__2_;
   wire DPATH_RF_MEMORY_6__3_;
   wire DPATH_RF_MEMORY_6__4_;
   wire DPATH_RF_MEMORY_6__5_;
   wire DPATH_RF_MEMORY_6__6_;
   wire DPATH_RF_MEMORY_6__7_;
   wire DPATH_RF_MEMORY_6__8_;
   wire DPATH_RF_MEMORY_6__9_;
   wire DPATH_RF_MEMORY_6__10_;
   wire DPATH_RF_MEMORY_6__11_;
   wire DPATH_RF_MEMORY_6__12_;
   wire DPATH_RF_MEMORY_6__13_;
   wire DPATH_RF_MEMORY_6__14_;
   wire DPATH_RF_MEMORY_6__15_;
   wire DPATH_RF_MEMORY_6__16_;
   wire DPATH_RF_MEMORY_6__17_;
   wire DPATH_RF_MEMORY_6__18_;
   wire DPATH_RF_MEMORY_6__19_;
   wire DPATH_RF_MEMORY_6__20_;
   wire DPATH_RF_MEMORY_6__21_;
   wire DPATH_RF_MEMORY_6__22_;
   wire DPATH_RF_MEMORY_6__23_;
   wire DPATH_RF_MEMORY_6__24_;
   wire DPATH_RF_MEMORY_6__25_;
   wire DPATH_RF_MEMORY_6__26_;
   wire DPATH_RF_MEMORY_6__27_;
   wire DPATH_RF_MEMORY_6__28_;
   wire DPATH_RF_MEMORY_6__29_;
   wire DPATH_RF_MEMORY_6__30_;
   wire DPATH_RF_MEMORY_6__31_;
   wire DPATH_RF_MEMORY_7__0_;
   wire DPATH_RF_MEMORY_7__1_;
   wire DPATH_RF_MEMORY_7__2_;
   wire DPATH_RF_MEMORY_7__3_;
   wire DPATH_RF_MEMORY_7__4_;
   wire DPATH_RF_MEMORY_7__5_;
   wire DPATH_RF_MEMORY_7__6_;
   wire DPATH_RF_MEMORY_7__7_;
   wire DPATH_RF_MEMORY_7__8_;
   wire DPATH_RF_MEMORY_7__9_;
   wire DPATH_RF_MEMORY_7__10_;
   wire DPATH_RF_MEMORY_7__11_;
   wire DPATH_RF_MEMORY_7__12_;
   wire DPATH_RF_MEMORY_7__13_;
   wire DPATH_RF_MEMORY_7__14_;
   wire DPATH_RF_MEMORY_7__15_;
   wire DPATH_RF_MEMORY_7__16_;
   wire DPATH_RF_MEMORY_7__17_;
   wire DPATH_RF_MEMORY_7__18_;
   wire DPATH_RF_MEMORY_7__19_;
   wire DPATH_RF_MEMORY_7__20_;
   wire DPATH_RF_MEMORY_7__21_;
   wire DPATH_RF_MEMORY_7__22_;
   wire DPATH_RF_MEMORY_7__23_;
   wire DPATH_RF_MEMORY_7__24_;
   wire DPATH_RF_MEMORY_7__25_;
   wire DPATH_RF_MEMORY_7__26_;
   wire DPATH_RF_MEMORY_7__27_;
   wire DPATH_RF_MEMORY_7__28_;
   wire DPATH_RF_MEMORY_7__29_;
   wire DPATH_RF_MEMORY_7__30_;
   wire DPATH_RF_MEMORY_7__31_;
   wire DPATH_RF_MEMORY_8__0_;
   wire DPATH_RF_MEMORY_8__1_;
   wire DPATH_RF_MEMORY_8__2_;
   wire DPATH_RF_MEMORY_8__3_;
   wire DPATH_RF_MEMORY_8__4_;
   wire DPATH_RF_MEMORY_8__5_;
   wire DPATH_RF_MEMORY_8__6_;
   wire DPATH_RF_MEMORY_8__7_;
   wire DPATH_RF_MEMORY_8__8_;
   wire DPATH_RF_MEMORY_8__9_;
   wire DPATH_RF_MEMORY_8__10_;
   wire DPATH_RF_MEMORY_8__11_;
   wire DPATH_RF_MEMORY_8__12_;
   wire DPATH_RF_MEMORY_8__13_;
   wire DPATH_RF_MEMORY_8__14_;
   wire DPATH_RF_MEMORY_8__15_;
   wire DPATH_RF_MEMORY_8__16_;
   wire DPATH_RF_MEMORY_8__17_;
   wire DPATH_RF_MEMORY_8__18_;
   wire DPATH_RF_MEMORY_8__19_;
   wire DPATH_RF_MEMORY_8__20_;
   wire DPATH_RF_MEMORY_8__21_;
   wire DPATH_RF_MEMORY_8__22_;
   wire DPATH_RF_MEMORY_8__23_;
   wire DPATH_RF_MEMORY_8__24_;
   wire DPATH_RF_MEMORY_8__25_;
   wire DPATH_RF_MEMORY_8__26_;
   wire DPATH_RF_MEMORY_8__27_;
   wire DPATH_RF_MEMORY_8__28_;
   wire DPATH_RF_MEMORY_8__29_;
   wire DPATH_RF_MEMORY_8__30_;
   wire DPATH_RF_MEMORY_8__31_;
   wire DPATH_RF_MEMORY_9__0_;
   wire DPATH_RF_MEMORY_9__1_;
   wire DPATH_RF_MEMORY_9__2_;
   wire DPATH_RF_MEMORY_9__3_;
   wire DPATH_RF_MEMORY_9__4_;
   wire DPATH_RF_MEMORY_9__5_;
   wire DPATH_RF_MEMORY_9__6_;
   wire DPATH_RF_MEMORY_9__7_;
   wire DPATH_RF_MEMORY_9__8_;
   wire DPATH_RF_MEMORY_9__9_;
   wire DPATH_RF_MEMORY_9__10_;
   wire DPATH_RF_MEMORY_9__11_;
   wire DPATH_RF_MEMORY_9__12_;
   wire DPATH_RF_MEMORY_9__13_;
   wire DPATH_RF_MEMORY_9__14_;
   wire DPATH_RF_MEMORY_9__15_;
   wire DPATH_RF_MEMORY_9__16_;
   wire DPATH_RF_MEMORY_9__17_;
   wire DPATH_RF_MEMORY_9__18_;
   wire DPATH_RF_MEMORY_9__19_;
   wire DPATH_RF_MEMORY_9__20_;
   wire DPATH_RF_MEMORY_9__21_;
   wire DPATH_RF_MEMORY_9__22_;
   wire DPATH_RF_MEMORY_9__23_;
   wire DPATH_RF_MEMORY_9__24_;
   wire DPATH_RF_MEMORY_9__25_;
   wire DPATH_RF_MEMORY_9__26_;
   wire DPATH_RF_MEMORY_9__27_;
   wire DPATH_RF_MEMORY_9__28_;
   wire DPATH_RF_MEMORY_9__29_;
   wire DPATH_RF_MEMORY_9__30_;
   wire DPATH_RF_MEMORY_9__31_;
   wire DPATH_RF_MEMORY_10__0_;
   wire DPATH_RF_MEMORY_10__1_;
   wire DPATH_RF_MEMORY_10__2_;
   wire DPATH_RF_MEMORY_10__3_;
   wire DPATH_RF_MEMORY_10__4_;
   wire DPATH_RF_MEMORY_10__5_;
   wire DPATH_RF_MEMORY_10__6_;
   wire DPATH_RF_MEMORY_10__7_;
   wire DPATH_RF_MEMORY_10__8_;
   wire DPATH_RF_MEMORY_10__9_;
   wire DPATH_RF_MEMORY_10__10_;
   wire DPATH_RF_MEMORY_10__11_;
   wire DPATH_RF_MEMORY_10__12_;
   wire DPATH_RF_MEMORY_10__13_;
   wire DPATH_RF_MEMORY_10__14_;
   wire DPATH_RF_MEMORY_10__15_;
   wire DPATH_RF_MEMORY_10__16_;
   wire DPATH_RF_MEMORY_10__17_;
   wire DPATH_RF_MEMORY_10__18_;
   wire DPATH_RF_MEMORY_10__19_;
   wire DPATH_RF_MEMORY_10__20_;
   wire DPATH_RF_MEMORY_10__21_;
   wire DPATH_RF_MEMORY_10__22_;
   wire DPATH_RF_MEMORY_10__23_;
   wire DPATH_RF_MEMORY_10__24_;
   wire DPATH_RF_MEMORY_10__25_;
   wire DPATH_RF_MEMORY_10__26_;
   wire DPATH_RF_MEMORY_10__27_;
   wire DPATH_RF_MEMORY_10__28_;
   wire DPATH_RF_MEMORY_10__29_;
   wire DPATH_RF_MEMORY_10__30_;
   wire DPATH_RF_MEMORY_10__31_;
   wire DPATH_RF_MEMORY_11__0_;
   wire DPATH_RF_MEMORY_11__1_;
   wire DPATH_RF_MEMORY_11__2_;
   wire DPATH_RF_MEMORY_11__3_;
   wire DPATH_RF_MEMORY_11__4_;
   wire DPATH_RF_MEMORY_11__5_;
   wire DPATH_RF_MEMORY_11__6_;
   wire DPATH_RF_MEMORY_11__7_;
   wire DPATH_RF_MEMORY_11__8_;
   wire DPATH_RF_MEMORY_11__9_;
   wire DPATH_RF_MEMORY_11__10_;
   wire DPATH_RF_MEMORY_11__11_;
   wire DPATH_RF_MEMORY_11__12_;
   wire DPATH_RF_MEMORY_11__13_;
   wire DPATH_RF_MEMORY_11__14_;
   wire DPATH_RF_MEMORY_11__15_;
   wire DPATH_RF_MEMORY_11__16_;
   wire DPATH_RF_MEMORY_11__17_;
   wire DPATH_RF_MEMORY_11__18_;
   wire DPATH_RF_MEMORY_11__19_;
   wire DPATH_RF_MEMORY_11__20_;
   wire DPATH_RF_MEMORY_11__21_;
   wire DPATH_RF_MEMORY_11__22_;
   wire DPATH_RF_MEMORY_11__23_;
   wire DPATH_RF_MEMORY_11__24_;
   wire DPATH_RF_MEMORY_11__25_;
   wire DPATH_RF_MEMORY_11__26_;
   wire DPATH_RF_MEMORY_11__27_;
   wire DPATH_RF_MEMORY_11__28_;
   wire DPATH_RF_MEMORY_11__29_;
   wire DPATH_RF_MEMORY_11__30_;
   wire DPATH_RF_MEMORY_11__31_;
   wire DPATH_RF_MEMORY_12__0_;
   wire DPATH_RF_MEMORY_12__1_;
   wire DPATH_RF_MEMORY_12__2_;
   wire DPATH_RF_MEMORY_12__3_;
   wire DPATH_RF_MEMORY_12__4_;
   wire DPATH_RF_MEMORY_12__5_;
   wire DPATH_RF_MEMORY_12__6_;
   wire DPATH_RF_MEMORY_12__7_;
   wire DPATH_RF_MEMORY_12__8_;
   wire DPATH_RF_MEMORY_12__9_;
   wire DPATH_RF_MEMORY_12__10_;
   wire DPATH_RF_MEMORY_12__11_;
   wire DPATH_RF_MEMORY_12__12_;
   wire DPATH_RF_MEMORY_12__13_;
   wire DPATH_RF_MEMORY_12__14_;
   wire DPATH_RF_MEMORY_12__15_;
   wire DPATH_RF_MEMORY_12__16_;
   wire DPATH_RF_MEMORY_12__17_;
   wire DPATH_RF_MEMORY_12__18_;
   wire DPATH_RF_MEMORY_12__19_;
   wire DPATH_RF_MEMORY_12__20_;
   wire DPATH_RF_MEMORY_12__21_;
   wire DPATH_RF_MEMORY_12__22_;
   wire DPATH_RF_MEMORY_12__23_;
   wire DPATH_RF_MEMORY_12__24_;
   wire DPATH_RF_MEMORY_12__25_;
   wire DPATH_RF_MEMORY_12__26_;
   wire DPATH_RF_MEMORY_12__27_;
   wire DPATH_RF_MEMORY_12__28_;
   wire DPATH_RF_MEMORY_12__29_;
   wire DPATH_RF_MEMORY_12__30_;
   wire DPATH_RF_MEMORY_12__31_;
   wire DPATH_RF_MEMORY_13__0_;
   wire DPATH_RF_MEMORY_13__1_;
   wire DPATH_RF_MEMORY_13__2_;
   wire DPATH_RF_MEMORY_13__3_;
   wire DPATH_RF_MEMORY_13__4_;
   wire DPATH_RF_MEMORY_13__5_;
   wire DPATH_RF_MEMORY_13__6_;
   wire DPATH_RF_MEMORY_13__7_;
   wire DPATH_RF_MEMORY_13__8_;
   wire DPATH_RF_MEMORY_13__9_;
   wire DPATH_RF_MEMORY_13__10_;
   wire DPATH_RF_MEMORY_13__11_;
   wire DPATH_RF_MEMORY_13__12_;
   wire DPATH_RF_MEMORY_13__13_;
   wire DPATH_RF_MEMORY_13__14_;
   wire DPATH_RF_MEMORY_13__15_;
   wire DPATH_RF_MEMORY_13__16_;
   wire DPATH_RF_MEMORY_13__17_;
   wire DPATH_RF_MEMORY_13__18_;
   wire DPATH_RF_MEMORY_13__19_;
   wire DPATH_RF_MEMORY_13__20_;
   wire DPATH_RF_MEMORY_13__21_;
   wire DPATH_RF_MEMORY_13__22_;
   wire DPATH_RF_MEMORY_13__23_;
   wire DPATH_RF_MEMORY_13__24_;
   wire DPATH_RF_MEMORY_13__25_;
   wire DPATH_RF_MEMORY_13__26_;
   wire DPATH_RF_MEMORY_13__27_;
   wire DPATH_RF_MEMORY_13__28_;
   wire DPATH_RF_MEMORY_13__29_;
   wire DPATH_RF_MEMORY_13__30_;
   wire DPATH_RF_MEMORY_13__31_;
   wire DPATH_RF_MEMORY_14__0_;
   wire DPATH_RF_MEMORY_14__1_;
   wire DPATH_RF_MEMORY_14__2_;
   wire DPATH_RF_MEMORY_14__3_;
   wire DPATH_RF_MEMORY_14__4_;
   wire DPATH_RF_MEMORY_14__5_;
   wire DPATH_RF_MEMORY_14__6_;
   wire DPATH_RF_MEMORY_14__7_;
   wire DPATH_RF_MEMORY_14__8_;
   wire DPATH_RF_MEMORY_14__9_;
   wire DPATH_RF_MEMORY_14__10_;
   wire DPATH_RF_MEMORY_14__11_;
   wire DPATH_RF_MEMORY_14__12_;
   wire DPATH_RF_MEMORY_14__13_;
   wire DPATH_RF_MEMORY_14__14_;
   wire DPATH_RF_MEMORY_14__15_;
   wire DPATH_RF_MEMORY_14__16_;
   wire DPATH_RF_MEMORY_14__17_;
   wire DPATH_RF_MEMORY_14__18_;
   wire DPATH_RF_MEMORY_14__19_;
   wire DPATH_RF_MEMORY_14__20_;
   wire DPATH_RF_MEMORY_14__21_;
   wire DPATH_RF_MEMORY_14__22_;
   wire DPATH_RF_MEMORY_14__23_;
   wire DPATH_RF_MEMORY_14__24_;
   wire DPATH_RF_MEMORY_14__25_;
   wire DPATH_RF_MEMORY_14__26_;
   wire DPATH_RF_MEMORY_14__27_;
   wire DPATH_RF_MEMORY_14__28_;
   wire DPATH_RF_MEMORY_14__29_;
   wire DPATH_RF_MEMORY_14__30_;
   wire DPATH_RF_MEMORY_14__31_;
   wire DPATH_RF_MEMORY_15__0_;
   wire DPATH_RF_MEMORY_15__1_;
   wire DPATH_RF_MEMORY_15__2_;
   wire DPATH_RF_MEMORY_15__3_;
   wire DPATH_RF_MEMORY_15__4_;
   wire DPATH_RF_MEMORY_15__5_;
   wire DPATH_RF_MEMORY_15__6_;
   wire DPATH_RF_MEMORY_15__7_;
   wire DPATH_RF_MEMORY_15__8_;
   wire DPATH_RF_MEMORY_15__9_;
   wire DPATH_RF_MEMORY_15__10_;
   wire DPATH_RF_MEMORY_15__11_;
   wire DPATH_RF_MEMORY_15__12_;
   wire DPATH_RF_MEMORY_15__13_;
   wire DPATH_RF_MEMORY_15__14_;
   wire DPATH_RF_MEMORY_15__15_;
   wire DPATH_RF_MEMORY_15__16_;
   wire DPATH_RF_MEMORY_15__17_;
   wire DPATH_RF_MEMORY_15__18_;
   wire DPATH_RF_MEMORY_15__19_;
   wire DPATH_RF_MEMORY_15__20_;
   wire DPATH_RF_MEMORY_15__21_;
   wire DPATH_RF_MEMORY_15__22_;
   wire DPATH_RF_MEMORY_15__23_;
   wire DPATH_RF_MEMORY_15__24_;
   wire DPATH_RF_MEMORY_15__25_;
   wire DPATH_RF_MEMORY_15__26_;
   wire DPATH_RF_MEMORY_15__27_;
   wire DPATH_RF_MEMORY_15__28_;
   wire DPATH_RF_MEMORY_15__29_;
   wire DPATH_RF_MEMORY_15__30_;
   wire DPATH_RF_MEMORY_15__31_;
   wire DPATH_RF_MEMORY_16__0_;
   wire DPATH_RF_MEMORY_16__1_;
   wire DPATH_RF_MEMORY_16__2_;
   wire DPATH_RF_MEMORY_16__3_;
   wire DPATH_RF_MEMORY_16__4_;
   wire DPATH_RF_MEMORY_16__5_;
   wire DPATH_RF_MEMORY_16__6_;
   wire DPATH_RF_MEMORY_16__7_;
   wire DPATH_RF_MEMORY_16__8_;
   wire DPATH_RF_MEMORY_16__9_;
   wire DPATH_RF_MEMORY_16__10_;
   wire DPATH_RF_MEMORY_16__11_;
   wire DPATH_RF_MEMORY_16__12_;
   wire DPATH_RF_MEMORY_16__13_;
   wire DPATH_RF_MEMORY_16__14_;
   wire DPATH_RF_MEMORY_16__15_;
   wire DPATH_RF_MEMORY_16__16_;
   wire DPATH_RF_MEMORY_16__17_;
   wire DPATH_RF_MEMORY_16__18_;
   wire DPATH_RF_MEMORY_16__19_;
   wire DPATH_RF_MEMORY_16__20_;
   wire DPATH_RF_MEMORY_16__21_;
   wire DPATH_RF_MEMORY_16__22_;
   wire DPATH_RF_MEMORY_16__23_;
   wire DPATH_RF_MEMORY_16__24_;
   wire DPATH_RF_MEMORY_16__25_;
   wire DPATH_RF_MEMORY_16__26_;
   wire DPATH_RF_MEMORY_16__27_;
   wire DPATH_RF_MEMORY_16__28_;
   wire DPATH_RF_MEMORY_16__29_;
   wire DPATH_RF_MEMORY_16__30_;
   wire DPATH_RF_MEMORY_16__31_;
   wire DPATH_RF_MEMORY_17__0_;
   wire DPATH_RF_MEMORY_17__1_;
   wire DPATH_RF_MEMORY_17__2_;
   wire DPATH_RF_MEMORY_17__3_;
   wire DPATH_RF_MEMORY_17__4_;
   wire DPATH_RF_MEMORY_17__5_;
   wire DPATH_RF_MEMORY_17__6_;
   wire DPATH_RF_MEMORY_17__7_;
   wire DPATH_RF_MEMORY_17__8_;
   wire DPATH_RF_MEMORY_17__9_;
   wire DPATH_RF_MEMORY_17__10_;
   wire DPATH_RF_MEMORY_17__11_;
   wire DPATH_RF_MEMORY_17__12_;
   wire DPATH_RF_MEMORY_17__13_;
   wire DPATH_RF_MEMORY_17__14_;
   wire DPATH_RF_MEMORY_17__15_;
   wire DPATH_RF_MEMORY_17__16_;
   wire DPATH_RF_MEMORY_17__17_;
   wire DPATH_RF_MEMORY_17__18_;
   wire DPATH_RF_MEMORY_17__19_;
   wire DPATH_RF_MEMORY_17__20_;
   wire DPATH_RF_MEMORY_17__21_;
   wire DPATH_RF_MEMORY_17__22_;
   wire DPATH_RF_MEMORY_17__23_;
   wire DPATH_RF_MEMORY_17__24_;
   wire DPATH_RF_MEMORY_17__25_;
   wire DPATH_RF_MEMORY_17__26_;
   wire DPATH_RF_MEMORY_17__27_;
   wire DPATH_RF_MEMORY_17__28_;
   wire DPATH_RF_MEMORY_17__29_;
   wire DPATH_RF_MEMORY_17__30_;
   wire DPATH_RF_MEMORY_17__31_;
   wire DPATH_RF_MEMORY_18__0_;
   wire DPATH_RF_MEMORY_18__1_;
   wire DPATH_RF_MEMORY_18__2_;
   wire DPATH_RF_MEMORY_18__3_;
   wire DPATH_RF_MEMORY_18__4_;
   wire DPATH_RF_MEMORY_18__5_;
   wire DPATH_RF_MEMORY_18__6_;
   wire DPATH_RF_MEMORY_18__7_;
   wire DPATH_RF_MEMORY_18__8_;
   wire DPATH_RF_MEMORY_18__9_;
   wire DPATH_RF_MEMORY_18__10_;
   wire DPATH_RF_MEMORY_18__11_;
   wire DPATH_RF_MEMORY_18__12_;
   wire DPATH_RF_MEMORY_18__13_;
   wire DPATH_RF_MEMORY_18__14_;
   wire DPATH_RF_MEMORY_18__15_;
   wire DPATH_RF_MEMORY_18__16_;
   wire DPATH_RF_MEMORY_18__17_;
   wire DPATH_RF_MEMORY_18__18_;
   wire DPATH_RF_MEMORY_18__19_;
   wire DPATH_RF_MEMORY_18__20_;
   wire DPATH_RF_MEMORY_18__21_;
   wire DPATH_RF_MEMORY_18__22_;
   wire DPATH_RF_MEMORY_18__23_;
   wire DPATH_RF_MEMORY_18__24_;
   wire DPATH_RF_MEMORY_18__25_;
   wire DPATH_RF_MEMORY_18__26_;
   wire DPATH_RF_MEMORY_18__27_;
   wire DPATH_RF_MEMORY_18__28_;
   wire DPATH_RF_MEMORY_18__29_;
   wire DPATH_RF_MEMORY_18__30_;
   wire DPATH_RF_MEMORY_18__31_;
   wire DPATH_RF_MEMORY_19__0_;
   wire DPATH_RF_MEMORY_19__1_;
   wire DPATH_RF_MEMORY_19__2_;
   wire DPATH_RF_MEMORY_19__3_;
   wire DPATH_RF_MEMORY_19__4_;
   wire DPATH_RF_MEMORY_19__5_;
   wire DPATH_RF_MEMORY_19__6_;
   wire DPATH_RF_MEMORY_19__7_;
   wire DPATH_RF_MEMORY_19__8_;
   wire DPATH_RF_MEMORY_19__9_;
   wire DPATH_RF_MEMORY_19__10_;
   wire DPATH_RF_MEMORY_19__11_;
   wire DPATH_RF_MEMORY_19__12_;
   wire DPATH_RF_MEMORY_19__13_;
   wire DPATH_RF_MEMORY_19__14_;
   wire DPATH_RF_MEMORY_19__15_;
   wire DPATH_RF_MEMORY_19__16_;
   wire DPATH_RF_MEMORY_19__17_;
   wire DPATH_RF_MEMORY_19__18_;
   wire DPATH_RF_MEMORY_19__19_;
   wire DPATH_RF_MEMORY_19__20_;
   wire DPATH_RF_MEMORY_19__21_;
   wire DPATH_RF_MEMORY_19__22_;
   wire DPATH_RF_MEMORY_19__23_;
   wire DPATH_RF_MEMORY_19__24_;
   wire DPATH_RF_MEMORY_19__25_;
   wire DPATH_RF_MEMORY_19__26_;
   wire DPATH_RF_MEMORY_19__27_;
   wire DPATH_RF_MEMORY_19__28_;
   wire DPATH_RF_MEMORY_19__29_;
   wire DPATH_RF_MEMORY_19__30_;
   wire DPATH_RF_MEMORY_19__31_;
   wire DPATH_RF_MEMORY_20__0_;
   wire DPATH_RF_MEMORY_20__1_;
   wire DPATH_RF_MEMORY_20__2_;
   wire DPATH_RF_MEMORY_20__3_;
   wire DPATH_RF_MEMORY_20__4_;
   wire DPATH_RF_MEMORY_20__5_;
   wire DPATH_RF_MEMORY_20__6_;
   wire DPATH_RF_MEMORY_20__7_;
   wire DPATH_RF_MEMORY_20__8_;
   wire DPATH_RF_MEMORY_20__9_;
   wire DPATH_RF_MEMORY_20__10_;
   wire DPATH_RF_MEMORY_20__11_;
   wire DPATH_RF_MEMORY_20__12_;
   wire DPATH_RF_MEMORY_20__13_;
   wire DPATH_RF_MEMORY_20__14_;
   wire DPATH_RF_MEMORY_20__15_;
   wire DPATH_RF_MEMORY_20__16_;
   wire DPATH_RF_MEMORY_20__17_;
   wire DPATH_RF_MEMORY_20__18_;
   wire DPATH_RF_MEMORY_20__19_;
   wire DPATH_RF_MEMORY_20__20_;
   wire DPATH_RF_MEMORY_20__21_;
   wire DPATH_RF_MEMORY_20__22_;
   wire DPATH_RF_MEMORY_20__23_;
   wire DPATH_RF_MEMORY_20__24_;
   wire DPATH_RF_MEMORY_20__25_;
   wire DPATH_RF_MEMORY_20__26_;
   wire DPATH_RF_MEMORY_20__27_;
   wire DPATH_RF_MEMORY_20__28_;
   wire DPATH_RF_MEMORY_20__29_;
   wire DPATH_RF_MEMORY_20__30_;
   wire DPATH_RF_MEMORY_20__31_;
   wire DPATH_RF_MEMORY_21__0_;
   wire DPATH_RF_MEMORY_21__1_;
   wire DPATH_RF_MEMORY_21__2_;
   wire DPATH_RF_MEMORY_21__3_;
   wire DPATH_RF_MEMORY_21__4_;
   wire DPATH_RF_MEMORY_21__5_;
   wire DPATH_RF_MEMORY_21__6_;
   wire DPATH_RF_MEMORY_21__7_;
   wire DPATH_RF_MEMORY_21__8_;
   wire DPATH_RF_MEMORY_21__9_;
   wire DPATH_RF_MEMORY_21__10_;
   wire DPATH_RF_MEMORY_21__11_;
   wire DPATH_RF_MEMORY_21__12_;
   wire DPATH_RF_MEMORY_21__13_;
   wire DPATH_RF_MEMORY_21__14_;
   wire DPATH_RF_MEMORY_21__15_;
   wire DPATH_RF_MEMORY_21__16_;
   wire DPATH_RF_MEMORY_21__17_;
   wire DPATH_RF_MEMORY_21__18_;
   wire DPATH_RF_MEMORY_21__19_;
   wire DPATH_RF_MEMORY_21__20_;
   wire DPATH_RF_MEMORY_21__21_;
   wire DPATH_RF_MEMORY_21__22_;
   wire DPATH_RF_MEMORY_21__23_;
   wire DPATH_RF_MEMORY_21__24_;
   wire DPATH_RF_MEMORY_21__25_;
   wire DPATH_RF_MEMORY_21__26_;
   wire DPATH_RF_MEMORY_21__27_;
   wire DPATH_RF_MEMORY_21__28_;
   wire DPATH_RF_MEMORY_21__29_;
   wire DPATH_RF_MEMORY_21__30_;
   wire DPATH_RF_MEMORY_21__31_;
   wire DPATH_RF_MEMORY_22__0_;
   wire DPATH_RF_MEMORY_22__1_;
   wire DPATH_RF_MEMORY_22__2_;
   wire DPATH_RF_MEMORY_22__3_;
   wire DPATH_RF_MEMORY_22__4_;
   wire DPATH_RF_MEMORY_22__5_;
   wire DPATH_RF_MEMORY_22__6_;
   wire DPATH_RF_MEMORY_22__7_;
   wire DPATH_RF_MEMORY_22__8_;
   wire DPATH_RF_MEMORY_22__9_;
   wire DPATH_RF_MEMORY_22__10_;
   wire DPATH_RF_MEMORY_22__11_;
   wire DPATH_RF_MEMORY_22__12_;
   wire DPATH_RF_MEMORY_22__13_;
   wire DPATH_RF_MEMORY_22__14_;
   wire DPATH_RF_MEMORY_22__15_;
   wire DPATH_RF_MEMORY_22__16_;
   wire DPATH_RF_MEMORY_22__17_;
   wire DPATH_RF_MEMORY_22__18_;
   wire DPATH_RF_MEMORY_22__19_;
   wire DPATH_RF_MEMORY_22__20_;
   wire DPATH_RF_MEMORY_22__21_;
   wire DPATH_RF_MEMORY_22__22_;
   wire DPATH_RF_MEMORY_22__23_;
   wire DPATH_RF_MEMORY_22__24_;
   wire DPATH_RF_MEMORY_22__25_;
   wire DPATH_RF_MEMORY_22__26_;
   wire DPATH_RF_MEMORY_22__27_;
   wire DPATH_RF_MEMORY_22__28_;
   wire DPATH_RF_MEMORY_22__29_;
   wire DPATH_RF_MEMORY_22__30_;
   wire DPATH_RF_MEMORY_22__31_;
   wire DPATH_RF_MEMORY_23__0_;
   wire DPATH_RF_MEMORY_23__1_;
   wire DPATH_RF_MEMORY_23__2_;
   wire DPATH_RF_MEMORY_23__3_;
   wire DPATH_RF_MEMORY_23__4_;
   wire DPATH_RF_MEMORY_23__5_;
   wire DPATH_RF_MEMORY_23__6_;
   wire DPATH_RF_MEMORY_23__7_;
   wire DPATH_RF_MEMORY_23__8_;
   wire DPATH_RF_MEMORY_23__9_;
   wire DPATH_RF_MEMORY_23__10_;
   wire DPATH_RF_MEMORY_23__11_;
   wire DPATH_RF_MEMORY_23__12_;
   wire DPATH_RF_MEMORY_23__13_;
   wire DPATH_RF_MEMORY_23__14_;
   wire DPATH_RF_MEMORY_23__15_;
   wire DPATH_RF_MEMORY_23__16_;
   wire DPATH_RF_MEMORY_23__17_;
   wire DPATH_RF_MEMORY_23__18_;
   wire DPATH_RF_MEMORY_23__19_;
   wire DPATH_RF_MEMORY_23__20_;
   wire DPATH_RF_MEMORY_23__21_;
   wire DPATH_RF_MEMORY_23__22_;
   wire DPATH_RF_MEMORY_23__23_;
   wire DPATH_RF_MEMORY_23__24_;
   wire DPATH_RF_MEMORY_23__25_;
   wire DPATH_RF_MEMORY_23__26_;
   wire DPATH_RF_MEMORY_23__27_;
   wire DPATH_RF_MEMORY_23__28_;
   wire DPATH_RF_MEMORY_23__29_;
   wire DPATH_RF_MEMORY_23__30_;
   wire DPATH_RF_MEMORY_23__31_;
   wire DPATH_RF_MEMORY_24__0_;
   wire DPATH_RF_MEMORY_24__1_;
   wire DPATH_RF_MEMORY_24__2_;
   wire DPATH_RF_MEMORY_24__3_;
   wire DPATH_RF_MEMORY_24__4_;
   wire DPATH_RF_MEMORY_24__5_;
   wire DPATH_RF_MEMORY_24__6_;
   wire DPATH_RF_MEMORY_24__7_;
   wire DPATH_RF_MEMORY_24__8_;
   wire DPATH_RF_MEMORY_24__9_;
   wire DPATH_RF_MEMORY_24__10_;
   wire DPATH_RF_MEMORY_24__11_;
   wire DPATH_RF_MEMORY_24__12_;
   wire DPATH_RF_MEMORY_24__13_;
   wire DPATH_RF_MEMORY_24__14_;
   wire DPATH_RF_MEMORY_24__15_;
   wire DPATH_RF_MEMORY_24__16_;
   wire DPATH_RF_MEMORY_24__17_;
   wire DPATH_RF_MEMORY_24__18_;
   wire DPATH_RF_MEMORY_24__19_;
   wire DPATH_RF_MEMORY_24__20_;
   wire DPATH_RF_MEMORY_24__21_;
   wire DPATH_RF_MEMORY_24__22_;
   wire DPATH_RF_MEMORY_24__23_;
   wire DPATH_RF_MEMORY_24__24_;
   wire DPATH_RF_MEMORY_24__25_;
   wire DPATH_RF_MEMORY_24__26_;
   wire DPATH_RF_MEMORY_24__27_;
   wire DPATH_RF_MEMORY_24__28_;
   wire DPATH_RF_MEMORY_24__29_;
   wire DPATH_RF_MEMORY_24__30_;
   wire DPATH_RF_MEMORY_24__31_;
   wire DPATH_RF_MEMORY_25__0_;
   wire DPATH_RF_MEMORY_25__1_;
   wire DPATH_RF_MEMORY_25__2_;
   wire DPATH_RF_MEMORY_25__3_;
   wire DPATH_RF_MEMORY_25__4_;
   wire DPATH_RF_MEMORY_25__5_;
   wire DPATH_RF_MEMORY_25__6_;
   wire DPATH_RF_MEMORY_25__7_;
   wire DPATH_RF_MEMORY_25__8_;
   wire DPATH_RF_MEMORY_25__9_;
   wire DPATH_RF_MEMORY_25__10_;
   wire DPATH_RF_MEMORY_25__11_;
   wire DPATH_RF_MEMORY_25__12_;
   wire DPATH_RF_MEMORY_25__13_;
   wire DPATH_RF_MEMORY_25__14_;
   wire DPATH_RF_MEMORY_25__15_;
   wire DPATH_RF_MEMORY_25__16_;
   wire DPATH_RF_MEMORY_25__17_;
   wire DPATH_RF_MEMORY_25__18_;
   wire DPATH_RF_MEMORY_25__19_;
   wire DPATH_RF_MEMORY_25__20_;
   wire DPATH_RF_MEMORY_25__21_;
   wire DPATH_RF_MEMORY_25__22_;
   wire DPATH_RF_MEMORY_25__23_;
   wire DPATH_RF_MEMORY_25__24_;
   wire DPATH_RF_MEMORY_25__25_;
   wire DPATH_RF_MEMORY_25__26_;
   wire DPATH_RF_MEMORY_25__27_;
   wire DPATH_RF_MEMORY_25__28_;
   wire DPATH_RF_MEMORY_25__29_;
   wire DPATH_RF_MEMORY_25__30_;
   wire DPATH_RF_MEMORY_25__31_;
   wire DPATH_RF_MEMORY_26__0_;
   wire DPATH_RF_MEMORY_26__1_;
   wire DPATH_RF_MEMORY_26__2_;
   wire DPATH_RF_MEMORY_26__3_;
   wire DPATH_RF_MEMORY_26__4_;
   wire DPATH_RF_MEMORY_26__5_;
   wire DPATH_RF_MEMORY_26__6_;
   wire DPATH_RF_MEMORY_26__7_;
   wire DPATH_RF_MEMORY_26__8_;
   wire DPATH_RF_MEMORY_26__9_;
   wire DPATH_RF_MEMORY_26__10_;
   wire DPATH_RF_MEMORY_26__11_;
   wire DPATH_RF_MEMORY_26__12_;
   wire DPATH_RF_MEMORY_26__13_;
   wire DPATH_RF_MEMORY_26__14_;
   wire DPATH_RF_MEMORY_26__15_;
   wire DPATH_RF_MEMORY_26__16_;
   wire DPATH_RF_MEMORY_26__17_;
   wire DPATH_RF_MEMORY_26__18_;
   wire DPATH_RF_MEMORY_26__19_;
   wire DPATH_RF_MEMORY_26__20_;
   wire DPATH_RF_MEMORY_26__21_;
   wire DPATH_RF_MEMORY_26__22_;
   wire DPATH_RF_MEMORY_26__23_;
   wire DPATH_RF_MEMORY_26__24_;
   wire DPATH_RF_MEMORY_26__25_;
   wire DPATH_RF_MEMORY_26__26_;
   wire DPATH_RF_MEMORY_26__27_;
   wire DPATH_RF_MEMORY_26__28_;
   wire DPATH_RF_MEMORY_26__29_;
   wire DPATH_RF_MEMORY_26__30_;
   wire DPATH_RF_MEMORY_26__31_;
   wire DPATH_RF_MEMORY_27__0_;
   wire DPATH_RF_MEMORY_27__1_;
   wire DPATH_RF_MEMORY_27__2_;
   wire DPATH_RF_MEMORY_27__3_;
   wire DPATH_RF_MEMORY_27__4_;
   wire DPATH_RF_MEMORY_27__5_;
   wire DPATH_RF_MEMORY_27__6_;
   wire DPATH_RF_MEMORY_27__7_;
   wire DPATH_RF_MEMORY_27__8_;
   wire DPATH_RF_MEMORY_27__9_;
   wire DPATH_RF_MEMORY_27__10_;
   wire DPATH_RF_MEMORY_27__11_;
   wire DPATH_RF_MEMORY_27__12_;
   wire DPATH_RF_MEMORY_27__13_;
   wire DPATH_RF_MEMORY_27__14_;
   wire DPATH_RF_MEMORY_27__15_;
   wire DPATH_RF_MEMORY_27__16_;
   wire DPATH_RF_MEMORY_27__17_;
   wire DPATH_RF_MEMORY_27__18_;
   wire DPATH_RF_MEMORY_27__19_;
   wire DPATH_RF_MEMORY_27__20_;
   wire DPATH_RF_MEMORY_27__21_;
   wire DPATH_RF_MEMORY_27__22_;
   wire DPATH_RF_MEMORY_27__23_;
   wire DPATH_RF_MEMORY_27__24_;
   wire DPATH_RF_MEMORY_27__25_;
   wire DPATH_RF_MEMORY_27__26_;
   wire DPATH_RF_MEMORY_27__27_;
   wire DPATH_RF_MEMORY_27__28_;
   wire DPATH_RF_MEMORY_27__29_;
   wire DPATH_RF_MEMORY_27__30_;
   wire DPATH_RF_MEMORY_27__31_;
   wire DPATH_RF_MEMORY_28__0_;
   wire DPATH_RF_MEMORY_28__1_;
   wire DPATH_RF_MEMORY_28__2_;
   wire DPATH_RF_MEMORY_28__3_;
   wire DPATH_RF_MEMORY_28__4_;
   wire DPATH_RF_MEMORY_28__5_;
   wire DPATH_RF_MEMORY_28__6_;
   wire DPATH_RF_MEMORY_28__7_;
   wire DPATH_RF_MEMORY_28__8_;
   wire DPATH_RF_MEMORY_28__9_;
   wire DPATH_RF_MEMORY_28__10_;
   wire DPATH_RF_MEMORY_28__11_;
   wire DPATH_RF_MEMORY_28__12_;
   wire DPATH_RF_MEMORY_28__13_;
   wire DPATH_RF_MEMORY_28__14_;
   wire DPATH_RF_MEMORY_28__15_;
   wire DPATH_RF_MEMORY_28__16_;
   wire DPATH_RF_MEMORY_28__17_;
   wire DPATH_RF_MEMORY_28__18_;
   wire DPATH_RF_MEMORY_28__19_;
   wire DPATH_RF_MEMORY_28__20_;
   wire DPATH_RF_MEMORY_28__21_;
   wire DPATH_RF_MEMORY_28__22_;
   wire DPATH_RF_MEMORY_28__23_;
   wire DPATH_RF_MEMORY_28__24_;
   wire DPATH_RF_MEMORY_28__25_;
   wire DPATH_RF_MEMORY_28__26_;
   wire DPATH_RF_MEMORY_28__27_;
   wire DPATH_RF_MEMORY_28__28_;
   wire DPATH_RF_MEMORY_28__29_;
   wire DPATH_RF_MEMORY_28__30_;
   wire DPATH_RF_MEMORY_28__31_;
   wire DPATH_RF_MEMORY_29__0_;
   wire DPATH_RF_MEMORY_29__1_;
   wire DPATH_RF_MEMORY_29__2_;
   wire DPATH_RF_MEMORY_29__3_;
   wire DPATH_RF_MEMORY_29__4_;
   wire DPATH_RF_MEMORY_29__5_;
   wire DPATH_RF_MEMORY_29__6_;
   wire DPATH_RF_MEMORY_29__7_;
   wire DPATH_RF_MEMORY_29__8_;
   wire DPATH_RF_MEMORY_29__9_;
   wire DPATH_RF_MEMORY_29__10_;
   wire DPATH_RF_MEMORY_29__11_;
   wire DPATH_RF_MEMORY_29__12_;
   wire DPATH_RF_MEMORY_29__13_;
   wire DPATH_RF_MEMORY_29__14_;
   wire DPATH_RF_MEMORY_29__15_;
   wire DPATH_RF_MEMORY_29__16_;
   wire DPATH_RF_MEMORY_29__17_;
   wire DPATH_RF_MEMORY_29__18_;
   wire DPATH_RF_MEMORY_29__19_;
   wire DPATH_RF_MEMORY_29__20_;
   wire DPATH_RF_MEMORY_29__21_;
   wire DPATH_RF_MEMORY_29__22_;
   wire DPATH_RF_MEMORY_29__23_;
   wire DPATH_RF_MEMORY_29__24_;
   wire DPATH_RF_MEMORY_29__25_;
   wire DPATH_RF_MEMORY_29__26_;
   wire DPATH_RF_MEMORY_29__27_;
   wire DPATH_RF_MEMORY_29__28_;
   wire DPATH_RF_MEMORY_29__29_;
   wire DPATH_RF_MEMORY_29__30_;
   wire DPATH_RF_MEMORY_29__31_;
   wire DPATH_RF_MEMORY_30__0_;
   wire DPATH_RF_MEMORY_30__1_;
   wire DPATH_RF_MEMORY_30__2_;
   wire DPATH_RF_MEMORY_30__3_;
   wire DPATH_RF_MEMORY_30__4_;
   wire DPATH_RF_MEMORY_30__5_;
   wire DPATH_RF_MEMORY_30__6_;
   wire DPATH_RF_MEMORY_30__7_;
   wire DPATH_RF_MEMORY_30__8_;
   wire DPATH_RF_MEMORY_30__9_;
   wire DPATH_RF_MEMORY_30__10_;
   wire DPATH_RF_MEMORY_30__11_;
   wire DPATH_RF_MEMORY_30__12_;
   wire DPATH_RF_MEMORY_30__13_;
   wire DPATH_RF_MEMORY_30__14_;
   wire DPATH_RF_MEMORY_30__15_;
   wire DPATH_RF_MEMORY_30__16_;
   wire DPATH_RF_MEMORY_30__17_;
   wire DPATH_RF_MEMORY_30__18_;
   wire DPATH_RF_MEMORY_30__19_;
   wire DPATH_RF_MEMORY_30__20_;
   wire DPATH_RF_MEMORY_30__21_;
   wire DPATH_RF_MEMORY_30__22_;
   wire DPATH_RF_MEMORY_30__23_;
   wire DPATH_RF_MEMORY_30__24_;
   wire DPATH_RF_MEMORY_30__25_;
   wire DPATH_RF_MEMORY_30__26_;
   wire DPATH_RF_MEMORY_30__27_;
   wire DPATH_RF_MEMORY_30__28_;
   wire DPATH_RF_MEMORY_30__29_;
   wire DPATH_RF_MEMORY_30__30_;
   wire DPATH_RF_MEMORY_30__31_;
   wire DPATH_RF_MEMORY_31__0_;
   wire DPATH_RF_MEMORY_31__1_;
   wire DPATH_RF_MEMORY_31__2_;
   wire DPATH_RF_MEMORY_31__3_;
   wire DPATH_RF_MEMORY_31__4_;
   wire DPATH_RF_MEMORY_31__5_;
   wire DPATH_RF_MEMORY_31__6_;
   wire DPATH_RF_MEMORY_31__7_;
   wire DPATH_RF_MEMORY_31__8_;
   wire DPATH_RF_MEMORY_31__9_;
   wire DPATH_RF_MEMORY_31__10_;
   wire DPATH_RF_MEMORY_31__11_;
   wire DPATH_RF_MEMORY_31__12_;
   wire DPATH_RF_MEMORY_31__13_;
   wire DPATH_RF_MEMORY_31__14_;
   wire DPATH_RF_MEMORY_31__15_;
   wire DPATH_RF_MEMORY_31__16_;
   wire DPATH_RF_MEMORY_31__17_;
   wire DPATH_RF_MEMORY_31__18_;
   wire DPATH_RF_MEMORY_31__19_;
   wire DPATH_RF_MEMORY_31__20_;
   wire DPATH_RF_MEMORY_31__21_;
   wire DPATH_RF_MEMORY_31__22_;
   wire DPATH_RF_MEMORY_31__23_;
   wire DPATH_RF_MEMORY_31__24_;
   wire DPATH_RF_MEMORY_31__25_;
   wire DPATH_RF_MEMORY_31__26_;
   wire DPATH_RF_MEMORY_31__27_;
   wire DPATH_RF_MEMORY_31__28_;
   wire DPATH_RF_MEMORY_31__29_;
   wire DPATH_RF_MEMORY_31__30_;
   wire DPATH_RF_MEMORY_31__31_;
   wire DPATH_addinc_ALU_add_381_20_n_1104;
   wire DPATH_addinc_ALU_add_381_20_n_1106;
   wire DPATH_addinc_ALU_add_381_20_n_1108;
   wire DPATH_addinc_ALU_add_381_20_n_1110;
   wire DPATH_addinc_ALU_add_381_20_n_1112;
   wire DPATH_addinc_ALU_add_381_20_n_1114;
   wire DPATH_addinc_ALU_add_381_20_n_1116;
   wire DPATH_addinc_ALU_add_381_20_n_1118;
   wire DPATH_addinc_ALU_add_381_20_n_1120;
   wire DPATH_addinc_ALU_add_381_20_n_1122;
   wire DPATH_addinc_ALU_add_381_20_n_1124;
   wire DPATH_addinc_ALU_add_381_20_n_1126;
   wire DPATH_addinc_ALU_add_381_20_n_1128;
   wire DPATH_addinc_ALU_add_381_20_n_1130;
   wire DPATH_addinc_ALU_add_381_20_n_1132;
   wire DPATH_addinc_ALU_add_381_20_n_1134;
   wire DPATH_addinc_ALU_add_381_20_n_1136;
   wire DPATH_addinc_ALU_add_381_20_n_1138;
   wire DPATH_addinc_ALU_add_381_20_n_1140;
   wire DPATH_addinc_ALU_add_381_20_n_1142;
   wire DPATH_addinc_ALU_add_381_20_n_1144;
   wire DPATH_addinc_ALU_add_381_20_n_1146;
   wire DPATH_addinc_ALU_add_381_20_n_1148;
   wire DPATH_addinc_ALU_add_381_20_n_1150;
   wire DPATH_addinc_ALU_add_381_20_n_1152;
   wire DPATH_addinc_ALU_add_381_20_n_1154;
   wire DPATH_addinc_ALU_add_381_20_n_1156;
   wire DPATH_addinc_ALU_add_381_20_n_1158;
   wire DPATH_addinc_ALU_add_381_20_n_1160;
   wire DPATH_addinc_ALU_add_381_20_n_1162;
   wire DPATH_addinc_ALU_add_381_20_n_1165;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_0;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_1;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_2;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_3;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_4;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_5;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_6;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_7;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_8;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_9;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_10;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_11;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_12;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_13;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_14;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_15;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_16;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_17;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_18;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_19;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_20;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_21;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_22;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_23;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_24;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_25;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_26;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_27;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_28;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_29;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_30;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_31;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_32;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_33;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_34;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_35;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_36;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_37;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_38;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_39;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_40;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_41;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_42;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_43;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_44;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_45;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_46;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_47;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_48;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_49;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_50;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_51;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_52;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_53;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_54;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_55;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_56;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_57;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_58;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_59;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_60;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_61;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_62;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_63;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_64;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_65;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_66;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_67;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_68;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_69;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_70;
   wire DPATH_csa_tree_ALU_eq_397_21_groupi_n_71;
   wire DPATH_n_2384;
   wire DPATH_n_2385;
   wire DPATH_n_2386;
   wire DPATH_n_2387;
   wire DPATH_n_2388;
   wire DPATH_n_2389;
   wire DPATH_n_2390;
   wire DPATH_n_2391;
   wire DPATH_n_2392;
   wire DPATH_n_2393;
   wire DPATH_n_2394;
   wire DPATH_n_2395;
   wire DPATH_n_2396;
   wire DPATH_n_2397;
   wire DPATH_n_2398;
   wire DPATH_n_2399;
   wire DPATH_n_2400;
   wire DPATH_n_2401;
   wire DPATH_n_2402;
   wire DPATH_n_2403;
   wire DPATH_n_2404;
   wire DPATH_n_2405;
   wire DPATH_n_2406;
   wire DPATH_n_2407;
   wire DPATH_n_2408;
   wire DPATH_n_2409;
   wire DPATH_n_2410;
   wire DPATH_n_2411;
   wire DPATH_n_2412;
   wire DPATH_n_2413;
   wire DPATH_n_2414;
   wire DPATH_n_2496;
   wire DPATH_n_2498;
   wire DPATH_n_2500;
   wire DPATH_n_2502;
   wire DPATH_n_2504;
   wire DPATH_n_2506;
   wire DPATH_n_2508;
   wire DPATH_n_2510;
   wire DPATH_n_2512;
   wire DPATH_n_2514;
   wire DPATH_n_2516;
   wire DPATH_n_2518;
   wire DPATH_n_2520;
   wire DPATH_n_2522;
   wire DPATH_n_2524;
   wire DPATH_n_2526;
   wire DPATH_n_2528;
   wire DPATH_n_2530;
   wire DPATH_n_2532;
   wire DPATH_n_2534;
   wire DPATH_n_2536;
   wire DPATH_n_2538;
   wire DPATH_n_2540;
   wire DPATH_n_2542;
   wire DPATH_n_2544;
   wire DPATH_n_2546;
   wire DPATH_n_2548;
   wire DPATH_n_2550;
   wire DPATH_n_2552;
   wire DPATH_n_2554;
   wire DPATH_n_2556;
   wire DPATH_n_2567;
   wire DPATH_n_2568;
   wire DPATH_n_2569;
   wire DPATH_n_2570;
   wire DPATH_n_2571;
   wire DPATH_n_2572;
   wire DPATH_n_2573;
   wire DPATH_n_2574;
   wire DPATH_n_2575;
   wire DPATH_n_2576;
   wire DPATH_n_2577;
   wire DPATH_n_2578;
   wire DPATH_n_2579;
   wire DPATH_n_2580;
   wire DPATH_n_2581;
   wire DPATH_n_2582;
   wire DPATH_n_2583;
   wire DPATH_n_2584;
   wire DPATH_n_2585;
   wire DPATH_n_2586;
   wire DPATH_n_2587;
   wire DPATH_n_2588;
   wire DPATH_n_2589;
   wire DPATH_n_2590;
   wire DPATH_n_2591;
   wire DPATH_n_2592;
   wire DPATH_n_2593;
   wire DPATH_n_2594;
   wire DPATH_n_2595;
   wire DPATH_n_2596;
   wire DPATH_n_2597;
   wire DPATH_n_2758;
   wire DPATH_n_2759;
   wire DPATH_n_2760;
   wire DPATH_n_2761;
   wire DPATH_n_2762;
   wire DPATH_n_2763;
   wire DPATH_n_2764;
   wire DPATH_n_2765;
   wire DPATH_n_2766;
   wire DPATH_n_2767;
   wire DPATH_n_2768;
   wire DPATH_n_2769;
   wire DPATH_n_2770;
   wire DPATH_n_2771;
   wire DPATH_n_2772;
   wire DPATH_n_2773;
   wire DPATH_n_2774;
   wire DPATH_n_2775;
   wire DPATH_n_2776;
   wire DPATH_n_2777;
   wire DPATH_n_2778;
   wire DPATH_n_2779;
   wire DPATH_n_2780;
   wire DPATH_n_2781;
   wire DPATH_n_2782;
   wire DPATH_n_2783;
   wire DPATH_n_2784;
   wire DPATH_n_2785;
   wire DPATH_n_2786;
   wire DPATH_n_2787;
   wire DPATH_n_2788;
   wire DPATH_n_2789;
   wire DPATH_n_2796;
   wire DPATH_n_2797;
   wire DPATH_n_2798;
   wire DPATH_n_2799;
   wire DPATH_n_2800;
   wire DPATH_n_2801;
   wire DPATH_n_2802;
   wire DPATH_n_2803;
   wire DPATH_n_2804;
   wire DPATH_n_2805;
   wire DPATH_n_2806;
   wire DPATH_n_2807;
   wire DPATH_n_2808;
   wire DPATH_n_2809;
   wire DPATH_n_2810;
   wire DPATH_n_2811;
   wire DPATH_n_2812;
   wire DPATH_n_2813;
   wire DPATH_n_2814;
   wire DPATH_n_2815;
   wire DPATH_n_2816;
   wire DPATH_n_2817;
   wire DPATH_n_2818;
   wire DPATH_n_2819;
   wire DPATH_n_2820;
   wire DPATH_n_2821;
   wire DPATH_n_2822;
   wire DPATH_n_2823;
   wire DPATH_n_2824;
   wire DPATH_n_2825;
   wire DPATH_n_2826;
   wire DPATH_n_2827;
   wire DPATH_n_2861;
   wire DPATH_n_2862;
   wire DPATH_n_2863;
   wire DPATH_n_2864;
   wire DPATH_n_2865;
   wire DPATH_n_2866;
   wire DPATH_n_2867;
   wire DPATH_n_2868;
   wire DPATH_n_2869;
   wire DPATH_n_2870;
   wire DPATH_n_2871;
   wire DPATH_n_2872;
   wire DPATH_n_2873;
   wire DPATH_n_2874;
   wire DPATH_n_2875;
   wire DPATH_n_2876;
   wire DPATH_n_2877;
   wire DPATH_n_2878;
   wire DPATH_n_2879;
   wire DPATH_n_2880;
   wire DPATH_n_2881;
   wire DPATH_n_2882;
   wire DPATH_n_2883;
   wire DPATH_n_2884;
   wire DPATH_n_2885;
   wire DPATH_n_2886;
   wire DPATH_n_2887;
   wire DPATH_n_2888;
   wire DPATH_n_2889;
   wire DPATH_n_2893;
   wire DPATH_n_2894;
   wire DPATH_n_2895;
   wire DPATH_n_2896;
   wire DPATH_n_2897;
   wire DPATH_n_2898;
   wire DPATH_n_2899;
   wire DPATH_n_2900;
   wire DPATH_n_2901;
   wire DPATH_n_2902;
   wire DPATH_n_2903;
   wire DPATH_n_2904;
   wire DPATH_n_2905;
   wire DPATH_n_2906;
   wire DPATH_n_2907;
   wire DPATH_n_2908;
   wire DPATH_n_2909;
   wire DPATH_n_2910;
   wire DPATH_n_2911;
   wire DPATH_n_2912;
   wire DPATH_n_2913;
   wire DPATH_n_2914;
   wire DPATH_n_2915;
   wire DPATH_n_2916;
   wire DPATH_n_2917;
   wire DPATH_n_2918;
   wire DPATH_n_2919;
   wire DPATH_n_2920;
   wire DPATH_n_2921;
   wire DPATH_n_2922;
   wire DPATH_n_2923;
   wire DPATH_n_5211;
   wire DPATH_n_5212;
   wire DPATH_n_5213;
   wire DPATH_n_5214;
   wire DPATH_n_5215;
   wire DPATH_n_5216;
   wire DPATH_n_5217;
   wire DPATH_n_5218;
   wire DPATH_n_5226;
   wire DPATH_n_5227;
   wire DPATH_n_5228;
   wire DPATH_n_5229;
   wire n_0;
   wire n_1;
   wire n_2;
   wire n_3;
   wire n_4;
   wire n_5;
   wire n_6;
   wire n_7;
   wire n_9;
   wire n_10;
   wire n_11;
   wire n_12;
   wire n_13;
   wire n_14;
   wire n_15;
   wire n_16;
   wire n_17;
   wire n_18;
   wire n_19;
   wire n_20;
   wire n_21;
   wire n_22;
   wire n_23;
   wire n_24;
   wire n_25;
   wire n_26;
   wire n_27;
   wire n_28;
   wire n_29;
   wire n_30;
   wire n_31;
   wire n_32;
   wire n_33;
   wire n_34;
   wire n_35;
   wire n_36;
   wire n_37;
   wire n_38;
   wire n_39;
   wire n_40;
   wire n_41;
   wire n_42;
   wire n_43;
   wire n_44;
   wire n_45;
   wire n_46;
   wire n_47;
   wire n_48;
   wire n_49;
   wire n_50;
   wire n_51;
   wire n_52;
   wire n_54;
   wire n_55;
   wire n_56;
   wire n_57;
   wire n_58;
   wire n_59;
   wire n_60;
   wire n_61;
   wire n_62;
   wire n_63;
   wire n_64;
   wire n_65;
   wire n_66;
   wire n_67;
   wire n_68;
   wire n_69;
   wire n_70;
   wire n_71;
   wire n_72;
   wire n_73;
   wire n_74;
   wire n_75;
   wire n_76;
   wire n_77;
   wire n_78;
   wire n_79;
   wire n_80;
   wire n_81;
   wire n_82;
   wire n_83;
   wire n_84;
   wire n_85;
   wire n_86;
   wire n_87;
   wire n_88;
   wire n_89;
   wire n_90;
   wire n_91;
   wire n_92;
   wire n_93;
   wire n_94;
   wire n_95;
   wire n_96;
   wire n_97;
   wire n_98;
   wire n_99;
   wire n_100;
   wire n_101;
   wire n_102;
   wire n_103;
   wire n_104;
   wire n_105;
   wire n_106;
   wire n_107;
   wire n_108;
   wire n_109;
   wire n_110;
   wire n_111;
   wire n_112;
   wire n_113;
   wire n_114;
   wire n_115;
   wire n_116;
   wire n_117;
   wire n_118;
   wire n_119;
   wire n_120;
   wire n_121;
   wire n_122;
   wire n_123;
   wire n_124;
   wire n_125;
   wire n_126;
   wire n_127;
   wire n_128;
   wire n_129;
   wire n_130;
   wire n_131;
   wire n_132;
   wire n_133;
   wire n_134;
   wire n_135;
   wire n_136;
   wire n_137;
   wire n_138;
   wire n_139;
   wire n_140;
   wire n_141;
   wire n_142;
   wire n_143;
   wire n_144;
   wire n_145;
   wire n_146;
   wire n_147;
   wire n_148;
   wire n_149;
   wire n_150;
   wire n_151;
   wire n_152;
   wire n_153;
   wire n_154;
   wire n_155;
   wire n_156;
   wire n_157;
   wire n_158;
   wire n_159;
   wire n_160;
   wire n_161;
   wire n_162;
   wire n_163;
   wire n_164;
   wire n_165;
   wire n_166;
   wire n_167;
   wire n_168;
   wire n_169;
   wire n_170;
   wire n_171;
   wire n_172;
   wire n_173;
   wire n_174;
   wire n_175;
   wire n_176;
   wire n_177;
   wire n_178;
   wire n_179;
   wire n_180;
   wire n_181;
   wire n_182;
   wire n_183;
   wire n_184;
   wire n_185;
   wire n_186;
   wire n_187;
   wire n_188;
   wire n_189;
   wire n_190;
   wire n_191;
   wire n_192;
   wire n_193;
   wire n_194;
   wire n_195;
   wire n_196;
   wire n_197;
   wire n_198;
   wire n_199;
   wire n_200;
   wire n_201;
   wire n_202;
   wire n_203;
   wire n_204;
   wire n_205;
   wire n_206;
   wire n_207;
   wire n_208;
   wire n_209;
   wire n_210;
   wire n_211;
   wire n_212;
   wire n_213;
   wire n_214;
   wire n_215;
   wire n_216;
   wire n_217;
   wire n_218;
   wire n_219;
   wire n_220;
   wire n_221;
   wire n_222;
   wire n_223;
   wire n_224;
   wire n_225;
   wire n_226;
   wire n_227;
   wire n_228;
   wire n_229;
   wire n_230;
   wire n_231;
   wire n_232;
   wire n_233;
   wire n_234;
   wire n_235;
   wire n_236;
   wire n_237;
   wire n_238;
   wire n_239;
   wire n_240;
   wire n_241;
   wire n_242;
   wire n_243;
   wire n_244;
   wire n_245;
   wire n_246;
   wire n_247;
   wire n_248;
   wire n_249;
   wire n_250;
   wire n_251;
   wire n_252;
   wire n_253;
   wire n_254;
   wire n_255;
   wire n_256;
   wire n_257;
   wire n_258;
   wire n_259;
   wire n_260;
   wire n_261;
   wire n_262;
   wire n_263;
   wire n_264;
   wire n_265;
   wire n_266;
   wire n_267;
   wire n_268;
   wire n_269;
   wire n_270;
   wire n_271;
   wire n_272;
   wire n_273;
   wire n_274;
   wire n_275;
   wire n_276;
   wire n_277;
   wire n_278;
   wire n_279;
   wire n_280;
   wire n_281;
   wire n_282;
   wire n_283;
   wire n_284;
   wire n_285;
   wire n_286;
   wire n_287;
   wire n_288;
   wire n_289;
   wire n_290;
   wire n_291;
   wire n_292;
   wire n_293;
   wire n_294;
   wire n_295;
   wire n_296;
   wire n_297;
   wire n_298;
   wire n_299;
   wire n_300;
   wire n_301;
   wire n_302;
   wire n_303;
   wire n_304;
   wire n_305;
   wire n_306;
   wire n_307;
   wire n_308;
   wire n_309;
   wire n_310;
   wire n_311;
   wire n_312;
   wire n_313;
   wire n_314;
   wire n_315;
   wire n_316;
   wire n_317;
   wire n_318;
   wire n_319;
   wire n_320;
   wire n_321;
   wire n_322;
   wire n_323;
   wire n_324;
   wire n_325;
   wire n_326;
   wire n_327;
   wire n_328;
   wire n_329;
   wire n_330;
   wire n_331;
   wire n_332;
   wire n_333;
   wire n_334;
   wire n_335;
   wire n_336;
   wire n_337;
   wire n_338;
   wire n_339;
   wire n_340;
   wire n_341;
   wire n_342;
   wire n_343;
   wire n_344;
   wire n_345;
   wire n_346;
   wire n_347;
   wire n_348;
   wire n_349;
   wire n_350;
   wire n_351;
   wire n_352;
   wire n_353;
   wire n_354;
   wire n_355;
   wire n_356;
   wire n_357;
   wire n_358;
   wire n_359;
   wire n_360;
   wire n_361;
   wire n_362;
   wire n_363;
   wire n_364;
   wire n_365;
   wire n_366;
   wire n_367;
   wire n_368;
   wire n_369;
   wire n_370;
   wire n_371;
   wire n_372;
   wire n_373;
   wire n_374;
   wire n_375;
   wire n_376;
   wire n_377;
   wire n_378;
   wire n_379;
   wire n_380;
   wire n_381;
   wire n_382;
   wire n_383;
   wire n_384;
   wire n_385;
   wire n_386;
   wire n_387;
   wire n_388;
   wire n_389;
   wire n_390;
   wire n_391;
   wire n_392;
   wire n_393;
   wire n_394;
   wire n_395;
   wire n_396;
   wire n_397;
   wire n_398;
   wire n_399;
   wire n_400;
   wire n_401;
   wire n_402;
   wire n_403;
   wire n_404;
   wire n_405;
   wire n_406;
   wire n_407;
   wire n_408;
   wire n_409;
   wire n_410;
   wire n_411;
   wire n_412;
   wire n_413;
   wire n_414;
   wire n_415;
   wire n_416;
   wire n_417;
   wire n_418;
   wire n_419;
   wire n_420;
   wire n_421;
   wire n_422;
   wire n_423;
   wire n_424;
   wire n_425;
   wire n_426;
   wire n_427;
   wire n_428;
   wire n_429;
   wire n_430;
   wire n_431;
   wire n_432;
   wire n_433;
   wire n_434;
   wire n_435;
   wire n_436;
   wire n_437;
   wire n_438;
   wire n_439;
   wire n_440;
   wire n_441;
   wire n_442;
   wire n_443;
   wire n_444;
   wire n_445;
   wire n_446;
   wire n_447;
   wire n_448;
   wire n_449;
   wire n_450;
   wire n_451;
   wire n_452;
   wire n_453;
   wire n_454;
   wire n_455;
   wire n_456;
   wire n_457;
   wire n_458;
   wire n_459;
   wire n_460;
   wire n_461;
   wire n_462;
   wire n_463;
   wire n_464;
   wire n_465;
   wire n_466;
   wire n_467;
   wire n_468;
   wire n_469;
   wire n_470;
   wire n_471;
   wire n_472;
   wire n_473;
   wire n_474;
   wire n_475;
   wire n_476;
   wire n_477;
   wire n_478;
   wire n_479;
   wire n_480;
   wire n_481;
   wire n_482;
   wire n_483;
   wire n_484;
   wire n_485;
   wire n_486;
   wire n_487;
   wire n_488;
   wire n_489;
   wire n_490;
   wire n_491;
   wire n_492;
   wire n_493;
   wire n_494;
   wire n_495;
   wire n_496;
   wire n_497;
   wire n_498;
   wire n_499;
   wire n_500;
   wire n_501;
   wire n_502;
   wire n_503;
   wire n_504;
   wire n_505;
   wire n_506;
   wire n_507;
   wire n_508;
   wire n_509;
   wire n_510;
   wire n_511;
   wire n_512;
   wire n_513;
   wire n_514;
   wire n_515;
   wire n_516;
   wire n_517;
   wire n_518;
   wire n_519;
   wire n_520;
   wire n_521;
   wire n_522;
   wire n_523;
   wire n_524;
   wire n_525;
   wire n_526;
   wire n_527;
   wire n_528;
   wire n_529;
   wire n_530;
   wire n_531;
   wire n_532;
   wire n_533;
   wire n_534;
   wire n_535;
   wire n_536;
   wire n_537;
   wire n_538;
   wire n_539;
   wire n_540;
   wire n_541;
   wire n_542;
   wire n_543;
   wire n_544;
   wire n_545;
   wire n_546;
   wire n_547;
   wire n_548;
   wire n_549;
   wire n_550;
   wire n_551;
   wire n_552;
   wire n_553;
   wire n_554;
   wire n_555;
   wire n_556;
   wire n_557;
   wire n_558;
   wire n_559;
   wire n_560;
   wire n_561;
   wire n_562;
   wire n_563;
   wire n_564;
   wire n_565;
   wire n_566;
   wire n_567;
   wire n_568;
   wire n_569;
   wire n_570;
   wire n_571;
   wire n_572;
   wire n_573;
   wire n_574;
   wire n_575;
   wire n_576;
   wire n_577;
   wire n_578;
   wire n_579;
   wire n_580;
   wire n_581;
   wire n_582;
   wire n_583;
   wire n_584;
   wire n_585;
   wire n_586;
   wire n_587;
   wire n_588;
   wire n_589;
   wire n_590;
   wire n_591;
   wire n_592;
   wire n_593;
   wire n_594;
   wire n_595;
   wire n_596;
   wire n_597;
   wire n_598;
   wire n_599;
   wire n_600;
   wire n_601;
   wire n_602;
   wire n_603;
   wire n_604;
   wire n_605;
   wire n_606;
   wire n_607;
   wire n_608;
   wire n_609;
   wire n_610;
   wire n_611;
   wire n_612;
   wire n_613;
   wire n_614;
   wire n_615;
   wire n_616;
   wire n_617;
   wire n_618;
   wire n_619;
   wire n_620;
   wire n_621;
   wire n_622;
   wire n_623;
   wire n_624;
   wire n_625;
   wire n_626;
   wire n_627;
   wire n_628;
   wire n_629;
   wire n_630;
   wire n_631;
   wire n_632;
   wire n_633;
   wire n_634;
   wire n_635;
   wire n_636;
   wire n_637;
   wire n_638;
   wire n_639;
   wire n_640;
   wire n_641;
   wire n_642;
   wire n_643;
   wire n_644;
   wire n_645;
   wire n_646;
   wire n_647;
   wire n_648;
   wire n_649;
   wire n_650;
   wire n_651;
   wire n_652;
   wire n_653;
   wire n_654;
   wire n_655;
   wire n_656;
   wire n_657;
   wire n_658;
   wire n_659;
   wire n_660;
   wire n_661;
   wire n_662;
   wire n_663;
   wire n_664;
   wire n_665;
   wire n_666;
   wire n_667;
   wire n_668;
   wire n_669;
   wire n_670;
   wire n_671;
   wire n_672;
   wire n_673;
   wire n_674;
   wire n_675;
   wire n_676;
   wire n_677;
   wire n_678;
   wire n_679;
   wire n_680;
   wire n_681;
   wire n_682;
   wire n_683;
   wire n_684;
   wire n_685;
   wire n_686;
   wire n_687;
   wire n_688;
   wire n_689;
   wire n_690;
   wire n_691;
   wire n_692;
   wire n_693;
   wire n_694;
   wire n_695;
   wire n_696;
   wire n_697;
   wire n_698;
   wire n_699;
   wire n_700;
   wire n_701;
   wire n_702;
   wire n_703;
   wire n_704;
   wire n_705;
   wire n_706;
   wire n_707;
   wire n_708;
   wire n_709;
   wire n_710;
   wire n_711;
   wire n_712;
   wire n_713;
   wire n_714;
   wire n_715;
   wire n_716;
   wire n_717;
   wire n_718;
   wire n_719;
   wire n_720;
   wire n_721;
   wire n_722;
   wire n_723;
   wire n_724;
   wire n_725;
   wire n_726;
   wire n_727;
   wire n_728;
   wire n_729;
   wire n_730;
   wire n_731;
   wire n_732;
   wire n_733;
   wire n_734;
   wire n_735;
   wire n_736;
   wire n_737;
   wire n_738;
   wire n_739;
   wire n_740;
   wire n_741;
   wire n_742;
   wire n_743;
   wire n_744;
   wire n_745;
   wire n_746;
   wire n_747;
   wire n_748;
   wire n_749;
   wire n_750;
   wire n_751;
   wire n_752;
   wire n_753;
   wire n_754;
   wire n_755;
   wire n_756;
   wire n_757;
   wire n_758;
   wire n_759;
   wire n_760;
   wire n_761;
   wire n_762;
   wire n_763;
   wire n_764;
   wire n_765;
   wire n_766;
   wire n_767;
   wire n_768;
   wire n_769;
   wire n_770;
   wire n_771;
   wire n_772;
   wire n_773;
   wire n_774;
   wire n_775;
   wire n_776;
   wire n_777;
   wire n_778;
   wire n_779;
   wire n_780;
   wire n_781;
   wire n_782;
   wire n_783;
   wire n_784;
   wire n_785;
   wire n_786;
   wire n_787;
   wire n_788;
   wire n_789;
   wire n_790;
   wire n_791;
   wire n_792;
   wire n_793;
   wire n_794;
   wire n_795;
   wire n_796;
   wire n_797;
   wire n_798;
   wire n_799;
   wire n_800;
   wire n_801;
   wire n_802;
   wire n_803;
   wire n_804;
   wire n_805;
   wire n_806;
   wire n_807;
   wire n_808;
   wire n_809;
   wire n_810;
   wire n_811;
   wire n_812;
   wire n_813;
   wire n_814;
   wire n_815;
   wire n_816;
   wire n_817;
   wire n_818;
   wire n_819;
   wire n_820;
   wire n_821;
   wire n_822;
   wire n_823;
   wire n_824;
   wire n_825;
   wire n_826;
   wire n_827;
   wire n_828;
   wire n_829;
   wire n_830;
   wire n_831;
   wire n_832;
   wire n_833;
   wire n_834;
   wire n_835;
   wire n_836;
   wire n_837;
   wire n_838;
   wire n_839;
   wire n_840;
   wire n_841;
   wire n_842;
   wire n_843;
   wire n_844;
   wire n_845;
   wire n_846;
   wire n_847;
   wire n_848;
   wire n_849;
   wire n_850;
   wire n_851;
   wire n_852;
   wire n_853;
   wire n_854;
   wire n_855;
   wire n_856;
   wire n_857;
   wire n_858;
   wire n_859;
   wire n_860;
   wire n_861;
   wire n_862;
   wire n_863;
   wire n_864;
   wire n_865;
   wire n_866;
   wire n_867;
   wire n_868;
   wire n_869;
   wire n_870;
   wire n_871;
   wire n_872;
   wire n_873;
   wire n_874;
   wire n_875;
   wire n_876;
   wire n_877;
   wire n_878;
   wire n_879;
   wire n_880;
   wire n_881;
   wire n_882;
   wire n_883;
   wire n_884;
   wire n_885;
   wire n_886;
   wire n_887;
   wire n_888;
   wire n_889;
   wire n_890;
   wire n_891;
   wire n_892;
   wire n_893;
   wire n_894;
   wire n_895;
   wire n_896;
   wire n_897;
   wire n_898;
   wire n_899;
   wire n_900;
   wire n_901;
   wire n_902;
   wire n_903;
   wire n_904;
   wire n_905;
   wire n_906;
   wire n_907;
   wire n_908;
   wire n_909;
   wire n_910;
   wire n_911;
   wire n_912;
   wire n_913;
   wire n_914;
   wire n_915;
   wire n_916;
   wire n_917;
   wire n_918;
   wire n_919;
   wire n_920;
   wire n_921;
   wire n_922;
   wire n_923;
   wire n_924;
   wire n_925;
   wire n_926;
   wire n_927;
   wire n_928;
   wire n_929;
   wire n_930;
   wire n_931;
   wire n_932;
   wire n_933;
   wire n_934;
   wire n_935;
   wire n_936;
   wire n_937;
   wire n_938;
   wire n_939;
   wire n_940;
   wire n_941;
   wire n_942;
   wire n_943;
   wire n_944;
   wire n_945;
   wire n_946;
   wire n_947;
   wire n_948;
   wire n_949;
   wire n_950;
   wire n_951;
   wire n_952;
   wire n_953;
   wire n_954;
   wire n_955;
   wire n_956;
   wire n_957;
   wire n_958;
   wire n_959;
   wire n_960;
   wire n_961;
   wire n_962;
   wire n_963;
   wire n_964;
   wire n_965;
   wire n_966;
   wire n_967;
   wire n_968;
   wire n_969;
   wire n_970;
   wire n_971;
   wire n_972;
   wire n_973;
   wire n_974;
   wire n_975;
   wire n_976;
   wire n_977;
   wire n_978;
   wire n_979;
   wire n_980;
   wire n_981;
   wire n_982;
   wire n_983;
   wire n_984;
   wire n_985;
   wire n_986;
   wire n_987;
   wire n_988;
   wire n_989;
   wire n_990;
   wire n_991;
   wire n_992;
   wire n_993;
   wire n_994;
   wire n_995;
   wire n_996;
   wire n_997;
   wire n_998;
   wire n_999;
   wire n_1000;
   wire n_1001;
   wire n_1002;
   wire n_1003;
   wire n_1004;
   wire n_1005;
   wire n_1006;
   wire n_1007;
   wire n_1008;
   wire n_1009;
   wire n_1010;
   wire n_1011;
   wire n_1012;
   wire n_1013;
   wire n_1014;
   wire n_1015;
   wire n_1016;
   wire n_1017;
   wire n_1018;
   wire n_1019;
   wire n_1020;
   wire n_1021;
   wire n_1022;
   wire n_1023;
   wire n_1024;
   wire n_1025;
   wire n_1026;
   wire n_1027;
   wire n_1028;
   wire n_1029;
   wire n_1030;
   wire n_1031;
   wire n_1032;
   wire n_1033;
   wire n_1034;
   wire n_1035;
   wire n_1036;
   wire n_1037;
   wire n_1038;
   wire n_1039;
   wire n_1040;
   wire n_1041;
   wire n_1042;
   wire n_1043;
   wire n_1044;
   wire n_1045;
   wire n_1046;
   wire n_1047;
   wire n_1048;
   wire n_1049;
   wire n_1050;
   wire n_1051;
   wire n_1052;
   wire n_1053;
   wire n_1054;
   wire n_1055;
   wire n_1056;
   wire n_1057;
   wire n_1058;
   wire n_1059;
   wire n_1060;
   wire n_1061;
   wire n_1062;
   wire n_1063;
   wire n_1064;
   wire n_1065;
   wire n_1066;
   wire n_1067;
   wire n_1068;
   wire n_1069;
   wire n_1070;
   wire n_1071;
   wire n_1072;
   wire n_1073;
   wire n_1074;
   wire n_1075;
   wire n_1076;
   wire n_1077;
   wire n_1078;
   wire n_1079;
   wire n_1080;
   wire n_1081;
   wire n_1082;
   wire n_1083;
   wire n_1084;
   wire n_1085;
   wire n_1086;
   wire n_1087;
   wire n_1088;
   wire n_1089;
   wire n_1090;
   wire n_1091;
   wire n_1092;
   wire n_1093;
   wire n_1094;
   wire n_1095;
   wire n_1096;
   wire n_1097;
   wire n_1098;
   wire n_1099;
   wire n_1100;
   wire n_1101;
   wire n_1102;
   wire n_1103;
   wire n_1104;
   wire n_1105;
   wire n_1106;
   wire n_1107;
   wire n_1108;
   wire n_1109;
   wire n_1110;
   wire n_1111;
   wire n_1112;
   wire n_1113;
   wire n_1114;
   wire n_1115;
   wire n_1116;
   wire n_1117;
   wire n_1118;
   wire n_1119;
   wire n_1120;
   wire n_1121;
   wire n_1122;
   wire n_1123;
   wire n_1124;
   wire n_1125;
   wire n_1126;
   wire n_1127;
   wire n_1128;
   wire n_1129;
   wire n_1130;
   wire n_1131;
   wire n_1132;
   wire n_1133;
   wire n_1134;
   wire n_1135;
   wire n_1136;
   wire n_1137;
   wire n_1138;
   wire n_1139;
   wire n_1140;
   wire n_1141;
   wire n_1142;
   wire n_1143;
   wire n_1144;
   wire n_1145;
   wire n_1146;
   wire n_1147;
   wire n_1148;
   wire n_1149;
   wire n_1150;
   wire n_1151;
   wire n_1152;
   wire n_1153;
   wire n_1154;
   wire n_1155;
   wire n_1156;
   wire n_1157;
   wire n_1158;
   wire n_1159;
   wire n_1160;
   wire n_1161;
   wire n_1162;
   wire n_1163;
   wire n_1164;
   wire n_1165;
   wire n_1166;
   wire n_1167;
   wire n_1168;
   wire n_1169;
   wire n_1170;
   wire n_1171;
   wire n_1172;
   wire n_1173;
   wire n_1174;
   wire n_1175;
   wire n_1176;
   wire n_1177;
   wire n_1178;
   wire n_1179;
   wire n_1180;
   wire n_1181;
   wire n_1182;
   wire n_1183;
   wire n_1184;
   wire n_1185;
   wire n_1186;
   wire n_1187;
   wire n_1188;
   wire n_1189;
   wire n_1190;
   wire n_1191;
   wire n_1192;
   wire n_1193;
   wire n_1194;
   wire n_1195;
   wire n_1196;
   wire n_1197;
   wire n_1198;
   wire n_1199;
   wire n_1200;
   wire n_1201;
   wire n_1202;
   wire n_1203;
   wire n_1204;
   wire n_1205;
   wire n_1206;
   wire n_1207;
   wire n_1208;
   wire n_1209;
   wire n_1210;
   wire n_1211;
   wire n_1212;
   wire n_1213;
   wire n_1214;
   wire n_1215;
   wire n_1216;
   wire n_1217;
   wire n_1218;
   wire n_1219;
   wire n_1220;
   wire n_1221;
   wire n_1222;
   wire n_1223;
   wire n_1224;
   wire n_1225;
   wire n_1226;
   wire n_1227;
   wire n_1228;
   wire n_1229;
   wire n_1230;
   wire n_1231;
   wire n_1232;
   wire n_1233;
   wire n_1234;
   wire n_1235;
   wire n_1236;
   wire n_1237;
   wire n_1238;
   wire n_1239;
   wire n_1240;
   wire n_1241;
   wire n_1242;
   wire n_1243;
   wire n_1244;
   wire n_1245;
   wire n_1246;
   wire n_1247;
   wire n_1248;
   wire n_1249;
   wire n_1250;
   wire n_1251;
   wire n_1252;
   wire n_1253;
   wire n_1254;
   wire n_1255;
   wire n_1256;
   wire n_1257;
   wire n_1258;
   wire n_1259;
   wire n_1260;
   wire n_1261;
   wire n_1262;
   wire n_1263;
   wire n_1264;
   wire n_1265;
   wire n_1266;
   wire n_1267;
   wire n_1268;
   wire n_1269;
   wire n_1270;
   wire n_1271;
   wire n_1272;
   wire n_1273;
   wire n_1274;
   wire n_1275;
   wire n_1276;
   wire n_1277;
   wire n_1278;
   wire n_1279;
   wire n_1280;
   wire n_1281;
   wire n_1282;
   wire n_1283;
   wire n_1284;
   wire n_1285;
   wire n_1286;
   wire n_1287;
   wire n_1288;
   wire n_1289;
   wire n_1290;
   wire n_1291;
   wire n_1292;
   wire n_1293;
   wire n_1294;
   wire n_1295;
   wire n_1296;
   wire n_1297;
   wire n_1298;
   wire n_1299;
   wire n_1300;
   wire n_1301;
   wire n_1302;
   wire n_1303;
   wire n_1304;
   wire n_1305;
   wire n_1306;
   wire n_1307;
   wire n_1308;
   wire n_1309;
   wire n_1310;
   wire n_1311;
   wire n_1312;
   wire n_1313;
   wire n_1314;
   wire n_1315;
   wire n_1316;
   wire n_1317;
   wire n_1318;
   wire n_1319;
   wire n_1320;
   wire n_1321;
   wire n_1322;
   wire n_1323;
   wire n_1324;
   wire n_1325;
   wire n_1326;
   wire n_1327;
   wire n_1328;
   wire n_1329;
   wire n_1330;
   wire n_1331;
   wire n_1332;
   wire n_1334;
   wire n_1335;
   wire n_1336;
   wire n_1337;
   wire n_1338;
   wire n_1339;
   wire n_1340;
   wire n_1341;
   wire n_1342;
   wire n_1343;
   wire n_1344;
   wire n_1345;
   wire n_1346;
   wire n_1347;
   wire n_1348;
   wire n_1349;
   wire n_1350;
   wire n_1351;
   wire n_1352;
   wire n_1353;
   wire n_1354;
   wire n_1355;
   wire n_1356;
   wire n_1357;
   wire n_1358;
   wire n_1360;
   wire n_1361;
   wire n_1362;
   wire n_1363;
   wire n_1364;
   wire n_1365;
   wire n_1366;
   wire n_1367;
   wire n_1368;
   wire n_1369;
   wire n_1371;
   wire n_1372;
   wire n_1373;
   wire n_1374;
   wire n_1375;
   wire n_1376;
   wire n_1377;
   wire n_1378;
   wire n_1379;
   wire n_1380;
   wire n_1381;
   wire n_1382;
   wire n_1383;
   wire n_1384;
   wire n_1385;
   wire n_1386;
   wire n_1387;
   wire n_1388;
   wire n_1389;
   wire n_1390;
   wire n_1391;
   wire n_1392;
   wire n_1393;
   wire n_1394;
   wire n_1395;
   wire n_1396;
   wire n_1397;
   wire n_1398;
   wire n_1399;
   wire n_1400;
   wire n_1401;
   wire n_1402;
   wire n_1403;
   wire n_1404;
   wire n_1405;
   wire n_1406;
   wire n_1407;
   wire n_1408;
   wire n_1409;
   wire n_1410;
   wire n_1411;
   wire n_1412;
   wire n_1413;
   wire n_1414;
   wire n_1415;
   wire n_1416;
   wire n_1417;
   wire n_1418;
   wire n_1419;
   wire n_1420;
   wire n_1421;
   wire n_1422;
   wire n_1423;
   wire n_1424;
   wire n_1425;
   wire n_1426;
   wire n_1427;
   wire n_1428;
   wire n_1429;
   wire n_1430;
   wire n_1431;
   wire n_1432;
   wire n_1433;
   wire n_1434;
   wire n_1435;
   wire n_1436;
   wire n_1437;
   wire n_1438;
   wire n_1439;
   wire n_1440;
   wire n_1441;
   wire n_1442;
   wire n_1443;
   wire n_1444;
   wire n_1445;
   wire n_1446;
   wire n_1447;
   wire n_1448;
   wire n_1449;
   wire n_1450;
   wire n_1451;
   wire n_1452;
   wire n_1453;
   wire n_1454;
   wire n_1455;
   wire n_1456;
   wire n_1457;
   wire n_1458;
   wire n_1459;
   wire n_1460;
   wire n_1461;
   wire n_1462;
   wire n_1463;
   wire n_1464;
   wire n_1465;
   wire n_1466;
   wire n_1468;
   wire n_1469;
   wire n_1470;
   wire n_1471;
   wire n_1472;
   wire n_1473;
   wire n_1474;
   wire n_1475;
   wire n_1476;
   wire n_1477;
   wire n_1478;
   wire n_1479;
   wire n_1480;
   wire n_1481;
   wire n_1482;
   wire n_1483;
   wire n_1484;
   wire n_1485;
   wire n_1486;
   wire n_1487;
   wire n_1488;
   wire n_1489;
   wire n_1490;
   wire n_1491;
   wire n_1492;
   wire n_1493;
   wire n_1494;
   wire n_1495;
   wire n_1496;
   wire n_1497;
   wire n_1498;
   wire n_1499;
   wire n_1500;
   wire n_1501;
   wire n_1502;
   wire n_1503;
   wire n_1504;
   wire n_1505;
   wire n_1506;
   wire n_1507;
   wire n_1508;
   wire n_1509;
   wire n_1510;
   wire n_1511;
   wire n_1512;
   wire n_1513;
   wire n_1514;
   wire n_1515;
   wire n_1516;
   wire n_1517;
   wire n_1518;
   wire n_1519;
   wire n_1520;
   wire n_1521;
   wire n_1522;
   wire n_1523;
   wire n_1524;
   wire n_1525;
   wire n_1526;
   wire n_1527;
   wire n_1528;
   wire n_1529;
   wire n_1530;
   wire n_1531;
   wire n_1532;
   wire n_1533;
   wire n_1534;
   wire n_1535;
   wire n_1536;
   wire n_1537;
   wire n_1538;
   wire n_1539;
   wire n_1540;
   wire n_1541;
   wire n_1542;
   wire n_1543;
   wire n_1544;
   wire n_1545;
   wire n_1546;
   wire n_1547;
   wire n_1548;
   wire n_1549;
   wire n_1550;
   wire n_1551;
   wire n_1552;
   wire n_1553;
   wire n_1554;
   wire n_1555;
   wire n_1556;
   wire n_1557;
   wire n_1558;
   wire n_1559;
   wire n_1560;
   wire n_1561;
   wire n_1562;
   wire n_1563;
   wire n_1564;
   wire n_1565;
   wire n_1566;
   wire n_1567;
   wire n_1568;
   wire n_1569;
   wire n_1570;
   wire n_1571;
   wire n_1572;
   wire n_1573;
   wire n_1574;
   wire n_1575;
   wire n_1576;
   wire n_1577;
   wire n_1578;
   wire n_1579;
   wire n_1580;
   wire n_1581;
   wire n_1582;
   wire n_1583;
   wire n_1584;
   wire n_1585;
   wire n_1586;
   wire n_1587;
   wire n_1588;
   wire n_1589;
   wire n_1590;
   wire n_1591;
   wire n_1592;
   wire n_1593;
   wire n_1594;
   wire n_1595;
   wire n_1596;
   wire n_1597;
   wire n_1598;
   wire n_1599;
   wire n_1600;
   wire n_1601;
   wire n_1602;
   wire n_1603;
   wire n_1604;
   wire n_1605;
   wire n_1606;
   wire n_1607;
   wire n_1608;
   wire n_1609;
   wire n_1610;
   wire n_1611;
   wire n_1612;
   wire n_1613;
   wire n_1614;
   wire n_1615;
   wire n_1616;
   wire n_1617;
   wire n_1618;
   wire n_1619;
   wire n_1620;
   wire n_1621;
   wire n_1622;
   wire n_1623;
   wire n_1624;
   wire n_1625;
   wire n_1626;
   wire n_1627;
   wire n_1628;
   wire n_1629;
   wire n_1630;
   wire n_1631;
   wire n_1632;
   wire n_1633;
   wire n_1634;
   wire n_1635;
   wire n_1636;
   wire n_1637;
   wire n_1638;
   wire n_1639;
   wire n_1640;
   wire n_1641;
   wire n_1642;
   wire n_1643;
   wire n_1644;
   wire n_1645;
   wire n_1646;
   wire n_1647;
   wire n_1648;
   wire n_1649;
   wire n_1650;
   wire n_1651;
   wire n_1652;
   wire n_1653;
   wire n_1654;
   wire n_1655;
   wire n_1656;
   wire n_1657;
   wire n_1658;
   wire n_1659;
   wire n_1660;
   wire n_1661;
   wire n_1662;
   wire n_1663;
   wire n_1664;
   wire n_1665;
   wire n_1666;
   wire n_1667;
   wire n_1668;
   wire n_1669;
   wire n_1670;
   wire n_1671;
   wire n_1672;
   wire n_1673;
   wire n_1674;
   wire n_1675;
   wire n_1676;
   wire n_1677;
   wire n_1678;
   wire n_1679;
   wire n_1680;
   wire n_1681;
   wire n_1682;
   wire n_1683;
   wire n_1684;
   wire n_1685;
   wire n_1686;
   wire n_1687;
   wire n_1688;
   wire n_1689;
   wire n_1690;
   wire n_1691;
   wire n_1692;
   wire n_1693;
   wire n_1694;
   wire n_1695;
   wire n_1696;
   wire n_1697;
   wire n_1698;
   wire n_1699;
   wire n_1700;
   wire n_1701;
   wire n_1702;
   wire n_1703;
   wire n_1704;
   wire n_1705;
   wire n_1706;
   wire n_1707;
   wire n_1708;
   wire n_1709;
   wire n_1710;
   wire n_1711;
   wire n_1712;
   wire n_1713;
   wire n_1714;
   wire n_1715;
   wire n_1716;
   wire n_1717;
   wire n_1718;
   wire n_1719;
   wire n_1720;
   wire n_1721;
   wire n_1722;
   wire n_1723;
   wire n_1724;
   wire n_1725;
   wire n_1726;
   wire n_1727;
   wire n_1728;
   wire n_1729;
   wire n_1730;
   wire n_1731;
   wire n_1732;
   wire n_1733;
   wire n_1734;
   wire n_1735;
   wire n_1736;
   wire n_1737;
   wire n_1738;
   wire n_1739;
   wire n_1740;
   wire n_1741;
   wire n_1742;
   wire n_1743;
   wire n_1744;
   wire n_1745;
   wire n_1746;
   wire n_1747;
   wire n_1748;
   wire n_1749;
   wire n_1750;
   wire n_1751;
   wire n_1752;
   wire n_1753;
   wire n_1754;
   wire n_1755;
   wire n_1756;
   wire n_1757;
   wire n_1758;
   wire n_1759;
   wire n_1760;
   wire n_1761;
   wire n_1762;
   wire n_1763;
   wire n_1764;
   wire n_1765;
   wire n_1766;
   wire n_1767;
   wire n_1768;
   wire n_1769;
   wire n_1770;
   wire n_1771;
   wire n_1772;
   wire n_1773;
   wire n_1774;
   wire n_1775;
   wire n_1776;
   wire n_1777;
   wire n_1778;
   wire n_1779;
   wire n_1780;
   wire n_1781;
   wire n_1782;
   wire n_1783;
   wire n_1784;
   wire n_1785;
   wire n_1786;
   wire n_1787;
   wire n_1788;
   wire n_1789;
   wire n_1790;
   wire n_1791;
   wire n_1792;
   wire n_1793;
   wire n_1794;
   wire n_1795;
   wire n_1796;
   wire n_1797;
   wire n_1798;
   wire n_1799;
   wire n_1800;
   wire n_1801;
   wire n_1802;
   wire n_1803;
   wire n_1804;
   wire n_1805;
   wire n_1806;
   wire n_1807;
   wire n_1808;
   wire n_1809;
   wire n_1810;
   wire n_1811;
   wire n_1812;
   wire n_1813;
   wire n_1814;
   wire n_1815;
   wire n_1816;
   wire n_1817;
   wire n_1818;
   wire n_1819;
   wire n_1820;
   wire n_1821;
   wire n_1822;
   wire n_1823;
   wire n_1824;
   wire n_1825;
   wire n_1826;
   wire n_1827;
   wire n_1828;
   wire n_1829;
   wire n_1830;
   wire n_1831;
   wire n_1832;
   wire n_1833;
   wire n_1834;
   wire n_1835;
   wire n_1836;
   wire n_1837;
   wire n_1838;
   wire n_1839;
   wire n_1840;
   wire n_1841;
   wire n_1842;
   wire n_1843;
   wire n_1844;
   wire n_1845;
   wire n_1846;
   wire n_1847;
   wire n_1848;
   wire n_1849;
   wire n_1850;
   wire n_1851;
   wire n_1852;
   wire n_1853;
   wire n_1854;
   wire n_1855;
   wire n_1856;
   wire n_1857;
   wire n_1858;
   wire n_1859;
   wire n_1860;
   wire n_1861;
   wire n_1862;
   wire n_1863;
   wire n_1864;
   wire n_1865;
   wire n_1866;
   wire n_1867;
   wire n_1868;
   wire n_1869;
   wire n_1870;
   wire n_1871;
   wire n_1872;
   wire n_1873;
   wire n_1874;
   wire n_1875;
   wire n_1876;
   wire n_1877;
   wire n_1878;
   wire n_1879;
   wire n_1880;
   wire n_1881;
   wire n_1882;
   wire n_1883;
   wire n_1884;
   wire n_1885;
   wire n_1886;
   wire n_1887;
   wire n_1888;
   wire n_1889;
   wire n_1890;
   wire n_1891;
   wire n_1892;
   wire n_1893;
   wire n_1894;
   wire n_1895;
   wire n_1896;
   wire n_1897;
   wire n_1898;
   wire n_1899;
   wire n_1900;
   wire n_1901;
   wire n_1902;
   wire n_1903;
   wire n_1904;
   wire n_1905;
   wire n_1906;
   wire n_1907;
   wire n_1908;
   wire n_1909;
   wire n_1910;
   wire n_1911;
   wire n_1912;
   wire n_1913;
   wire n_1914;
   wire n_1915;
   wire n_1916;
   wire n_1917;
   wire n_1918;
   wire n_1919;
   wire n_1920;
   wire n_1921;
   wire n_1922;
   wire n_1923;
   wire n_1924;
   wire n_1925;
   wire n_1926;
   wire n_1927;
   wire n_1928;
   wire n_1929;
   wire n_1930;
   wire n_1931;
   wire n_1932;
   wire n_1933;
   wire n_1934;
   wire n_1935;
   wire n_1936;
   wire n_1937;
   wire n_1938;
   wire n_1939;
   wire n_1940;
   wire n_1941;
   wire n_1942;
   wire n_1943;
   wire n_1944;
   wire n_1945;
   wire n_1946;
   wire n_1947;
   wire n_1948;
   wire n_1949;
   wire n_1950;
   wire n_1951;
   wire n_1952;
   wire n_1953;
   wire n_1954;
   wire n_1955;
   wire n_1956;
   wire n_1957;
   wire n_1958;
   wire n_1959;
   wire n_1960;
   wire n_1961;
   wire n_1962;
   wire n_1963;
   wire n_1964;
   wire n_1965;
   wire n_1966;
   wire n_1967;
   wire n_1968;
   wire n_1969;
   wire n_1970;
   wire n_1971;
   wire n_1972;
   wire n_1973;
   wire n_1974;
   wire n_1975;
   wire n_1976;
   wire n_1977;
   wire n_1978;
   wire n_1979;
   wire n_1980;
   wire n_1981;
   wire n_1982;
   wire n_1983;
   wire n_1984;
   wire n_1985;
   wire n_1986;
   wire n_1987;
   wire n_1988;
   wire n_1989;
   wire n_1990;
   wire n_1991;
   wire n_1992;
   wire n_1993;
   wire n_1994;
   wire n_1995;
   wire n_1996;
   wire n_1997;
   wire n_1998;
   wire n_1999;
   wire n_2000;
   wire n_2001;
   wire n_2002;
   wire n_2003;
   wire n_2004;
   wire n_2005;
   wire n_2006;
   wire n_2007;
   wire n_2008;
   wire n_2009;
   wire n_2010;
   wire n_2011;
   wire n_2012;
   wire n_2013;
   wire n_2014;
   wire n_2015;
   wire n_2016;
   wire n_2017;
   wire n_2018;
   wire n_2019;
   wire n_2020;
   wire n_2021;
   wire n_2022;
   wire n_2023;
   wire n_2024;
   wire n_2025;
   wire n_2026;
   wire n_2027;
   wire n_2028;
   wire n_2029;
   wire n_2030;
   wire n_2031;
   wire n_2032;
   wire n_2033;
   wire n_2034;
   wire n_2035;
   wire n_2036;
   wire n_2037;
   wire n_2038;
   wire n_2039;
   wire n_2040;
   wire n_2041;
   wire n_2042;
   wire n_2043;
   wire n_2044;
   wire n_2045;
   wire n_2046;
   wire n_2047;
   wire n_2048;
   wire n_2049;
   wire n_2050;
   wire n_2051;
   wire n_2052;
   wire n_2053;
   wire n_2054;
   wire n_2055;
   wire n_2056;
   wire n_2057;
   wire n_2058;
   wire n_2059;
   wire n_2060;
   wire n_2061;
   wire n_2062;
   wire n_2063;
   wire n_2064;
   wire n_2065;
   wire n_2066;
   wire n_2067;
   wire n_2068;
   wire n_2069;
   wire n_2070;
   wire n_2071;
   wire n_2072;
   wire n_2073;
   wire n_2074;
   wire n_2075;
   wire n_2076;
   wire n_2077;
   wire n_2078;
   wire n_2079;
   wire n_2080;
   wire n_2081;
   wire n_2082;
   wire n_2083;
   wire n_2084;
   wire n_2085;
   wire n_2086;
   wire n_2087;
   wire n_2088;
   wire n_2089;
   wire n_2090;
   wire n_2091;
   wire n_2092;
   wire n_2093;
   wire n_2094;
   wire n_2095;
   wire n_2096;
   wire n_2097;
   wire n_2098;
   wire n_2099;
   wire n_2100;
   wire n_2101;
   wire n_2102;
   wire n_2103;
   wire n_2104;
   wire n_2105;
   wire n_2106;
   wire n_2107;
   wire n_2108;
   wire n_2109;
   wire n_2110;
   wire n_2111;
   wire n_2112;
   wire n_2113;
   wire n_2114;
   wire n_2115;
   wire n_2116;
   wire n_2117;
   wire n_2118;
   wire n_2119;
   wire n_2120;
   wire n_2121;
   wire n_2122;
   wire n_2123;
   wire n_2124;
   wire n_2125;
   wire n_2126;
   wire n_2127;
   wire n_2128;
   wire n_2129;
   wire n_2130;
   wire n_2131;
   wire n_2132;
   wire n_2133;
   wire n_2134;
   wire n_2135;
   wire n_2136;
   wire n_2137;
   wire n_2138;
   wire n_2139;
   wire n_2140;
   wire n_2141;
   wire n_2142;
   wire n_2143;
   wire n_2144;
   wire n_2145;
   wire n_2146;
   wire n_2147;
   wire n_2148;
   wire n_2149;
   wire n_2150;
   wire n_2151;
   wire n_2152;
   wire n_2153;
   wire n_2154;
   wire n_2155;
   wire n_2156;
   wire n_2157;
   wire n_2158;
   wire n_2159;
   wire n_2160;
   wire n_2161;
   wire n_2162;
   wire n_2163;
   wire n_2164;
   wire n_2165;
   wire n_2166;
   wire n_2167;
   wire n_2168;
   wire n_2169;
   wire n_2170;
   wire n_2171;
   wire n_2172;
   wire n_2173;
   wire n_2174;
   wire n_2175;
   wire n_2176;
   wire n_2177;
   wire n_2178;
   wire n_2179;
   wire n_2180;
   wire n_2181;
   wire n_2182;
   wire n_2183;
   wire n_2184;
   wire n_2185;
   wire n_2186;
   wire n_2187;
   wire n_2188;
   wire n_2189;
   wire n_2190;
   wire n_2191;
   wire n_2192;
   wire n_2193;
   wire n_2194;
   wire n_2195;
   wire n_2196;
   wire n_2197;
   wire n_2198;
   wire n_2199;
   wire n_2200;
   wire n_2201;
   wire n_2202;
   wire n_2203;
   wire n_2204;
   wire n_2205;
   wire n_2206;
   wire n_2207;
   wire n_2209;
   wire n_2210;
   wire n_2211;
   wire n_2212;
   wire n_2213;
   wire n_2214;
   wire n_2215;
   wire n_2216;
   wire n_2217;
   wire n_2218;
   wire n_2219;
   wire n_2220;
   wire n_2221;
   wire n_2222;
   wire n_2223;
   wire n_2224;
   wire n_2225;
   wire n_2226;
   wire n_2227;
   wire n_2228;
   wire n_2229;
   wire n_2230;
   wire n_2231;
   wire n_2232;
   wire n_2233;
   wire n_2234;
   wire n_2235;
   wire n_2236;
   wire n_2237;
   wire n_2238;
   wire n_2239;
   wire n_2240;
   wire n_2241;
   wire n_2242;
   wire n_2243;
   wire n_2244;
   wire n_2245;
   wire n_2246;
   wire n_2247;
   wire n_2248;
   wire n_2249;
   wire n_2250;
   wire n_2251;
   wire n_2252;
   wire n_2253;
   wire n_2254;
   wire n_2255;
   wire n_2256;
   wire n_2257;
   wire n_2258;
   wire n_2259;
   wire n_2260;
   wire n_2261;
   wire n_2262;
   wire n_2263;
   wire n_2264;
   wire n_2265;
   wire n_2266;
   wire n_2267;
   wire n_2268;
   wire n_2269;
   wire n_2270;
   wire n_2271;
   wire n_2272;
   wire n_2273;
   wire n_2274;
   wire n_2275;
   wire n_2276;
   wire n_2277;
   wire n_2278;
   wire n_2279;
   wire n_2280;
   wire n_2281;
   wire n_2282;
   wire n_2283;
   wire n_2284;
   wire n_2285;
   wire n_2286;
   wire n_2287;
   wire n_2288;
   wire n_2289;
   wire n_2290;
   wire n_2291;
   wire n_2292;
   wire n_2293;
   wire n_2294;
   wire n_2295;
   wire n_2296;
   wire n_2297;
   wire n_2298;
   wire n_2299;
   wire n_2300;
   wire n_2301;
   wire n_2302;
   wire n_2303;
   wire n_2304;
   wire n_2305;
   wire n_2306;
   wire n_2307;
   wire n_2308;
   wire n_2309;
   wire n_2310;
   wire n_2311;
   wire n_2312;
   wire n_2313;
   wire n_2314;
   wire n_2315;
   wire n_2316;
   wire n_2317;
   wire n_2318;
   wire n_2319;
   wire n_2320;
   wire n_2321;
   wire n_2322;
   wire n_2323;
   wire n_2324;
   wire n_2325;
   wire n_2326;
   wire n_2327;
   wire n_2328;
   wire n_2329;
   wire n_2330;
   wire n_2331;
   wire n_2332;
   wire n_2333;
   wire n_2334;
   wire n_2335;
   wire n_2336;
   wire n_2337;
   wire n_2338;
   wire n_2339;
   wire n_2340;
   wire n_2341;
   wire n_2342;
   wire n_2343;
   wire n_2344;
   wire n_2345;
   wire n_2346;
   wire n_2347;
   wire n_2348;
   wire n_2349;
   wire n_2350;
   wire n_2351;
   wire n_2352;
   wire n_2353;
   wire n_2354;
   wire n_2355;
   wire n_2356;
   wire n_2357;
   wire n_2358;
   wire n_2359;
   wire n_2360;
   wire n_2361;
   wire n_2362;
   wire n_2363;
   wire n_2364;
   wire n_2365;
   wire n_2366;
   wire n_2367;
   wire n_2368;
   wire n_2369;
   wire n_2370;
   wire n_2371;
   wire n_2372;
   wire n_2373;
   wire n_2374;
   wire n_2375;
   wire n_2376;
   wire n_2377;
   wire n_2378;
   wire n_2379;
   wire n_2380;
   wire n_2381;
   wire n_2382;
   wire n_2383;
   wire n_2384;
   wire n_2385;
   wire n_2386;
   wire n_2387;
   wire n_2388;
   wire n_2389;
   wire n_2390;
   wire n_2391;
   wire n_2392;
   wire n_2393;
   wire n_2394;
   wire n_2395;
   wire n_2396;
   wire n_2397;
   wire n_2398;
   wire n_2399;
   wire n_2400;
   wire n_2401;
   wire n_2402;
   wire n_2403;
   wire n_2404;
   wire n_2405;
   wire n_2406;
   wire n_2407;
   wire n_2408;
   wire n_2409;
   wire n_2410;
   wire n_2411;
   wire n_2412;
   wire n_2413;
   wire n_2414;
   wire n_2415;
   wire n_2416;
   wire n_2417;
   wire n_2418;
   wire n_2419;
   wire n_2420;
   wire n_2421;
   wire n_2422;
   wire n_2423;
   wire n_2424;
   wire n_2425;
   wire n_2426;
   wire n_2427;
   wire n_2428;
   wire n_2429;
   wire n_2430;
   wire n_2431;
   wire n_2432;
   wire n_2433;
   wire n_2434;
   wire n_2435;
   wire n_2436;
   wire n_2437;
   wire n_2438;
   wire n_2439;
   wire n_2440;
   wire n_2441;
   wire n_2442;
   wire n_2443;
   wire n_2444;
   wire n_2445;
   wire n_2446;
   wire n_2447;
   wire n_2448;
   wire n_2449;
   wire n_2450;
   wire n_2451;
   wire n_2452;
   wire n_2453;
   wire n_2454;
   wire n_2455;
   wire n_2456;
   wire n_2457;
   wire n_2458;
   wire n_2459;
   wire n_2460;
   wire n_2461;
   wire n_2462;
   wire n_2463;
   wire n_2464;
   wire n_2465;
   wire n_2466;
   wire n_2467;
   wire n_2468;
   wire n_2469;
   wire n_2470;
   wire n_2471;
   wire n_2472;
   wire n_2473;
   wire n_2474;
   wire n_2475;
   wire n_2476;
   wire n_2477;
   wire n_2478;
   wire n_2479;
   wire n_2480;
   wire n_2481;
   wire n_2482;
   wire n_2483;
   wire n_2484;
   wire n_2485;
   wire n_2486;
   wire n_2487;
   wire n_2488;
   wire n_2489;
   wire n_2490;
   wire n_2491;
   wire n_2492;
   wire n_2493;
   wire n_2494;
   wire n_2495;
   wire n_2496;
   wire n_2497;
   wire n_2498;
   wire n_2499;
   wire n_2500;
   wire n_2501;
   wire n_2502;
   wire n_2503;
   wire n_2504;
   wire n_2505;
   wire n_2506;
   wire n_2507;
   wire n_2508;
   wire n_2509;
   wire n_2510;
   wire n_2511;
   wire n_2512;
   wire n_2513;
   wire n_2514;
   wire n_2515;
   wire n_2516;
   wire n_2517;
   wire n_2518;
   wire n_2519;
   wire n_2520;
   wire n_2521;
   wire n_2522;
   wire n_2523;
   wire n_2524;
   wire n_2525;
   wire n_2526;
   wire n_2527;
   wire n_2528;
   wire n_2529;
   wire n_2530;
   wire n_2531;
   wire n_2532;
   wire n_2533;
   wire n_2534;
   wire n_2535;
   wire n_2536;
   wire n_2537;
   wire n_2538;
   wire n_2539;
   wire n_2540;
   wire n_2541;
   wire n_2542;
   wire n_2543;
   wire n_2544;
   wire n_2545;
   wire n_2546;
   wire n_2547;
   wire n_2548;
   wire n_2549;
   wire n_2550;
   wire n_2551;
   wire n_2552;
   wire n_2553;
   wire n_2554;
   wire n_2555;
   wire n_2556;
   wire n_2557;
   wire n_2558;
   wire n_2559;
   wire n_2560;
   wire n_2561;
   wire n_2562;
   wire n_2563;
   wire n_2564;
   wire n_2565;
   wire n_2566;
   wire n_2567;
   wire n_2568;
   wire n_2569;
   wire n_2570;
   wire n_2571;
   wire n_2572;
   wire n_2573;
   wire n_2574;
   wire n_2575;
   wire n_2576;
   wire n_2577;
   wire n_2578;
   wire n_2579;
   wire n_2580;
   wire n_2581;
   wire n_2582;
   wire n_2583;
   wire n_2584;
   wire n_2585;
   wire n_2586;
   wire n_2587;
   wire n_2588;
   wire n_2589;
   wire n_2590;
   wire n_2591;
   wire n_2592;
   wire n_2593;
   wire n_2594;
   wire n_2595;
   wire n_2596;
   wire n_2597;
   wire n_2598;
   wire n_2599;
   wire n_2600;
   wire n_2601;
   wire n_2602;
   wire n_2603;
   wire n_2604;
   wire n_2605;
   wire n_2606;
   wire n_2607;
   wire n_2608;
   wire n_2609;
   wire n_2610;
   wire n_2611;
   wire n_2612;
   wire n_2613;
   wire n_2614;
   wire n_2615;
   wire n_2616;
   wire n_2617;
   wire n_2618;
   wire n_2619;
   wire n_2620;
   wire n_2621;
   wire n_2622;
   wire n_2623;
   wire n_2624;
   wire n_2625;
   wire n_2626;
   wire n_2627;
   wire n_2628;
   wire n_2629;
   wire n_2630;
   wire n_2631;
   wire n_2632;
   wire n_2633;
   wire n_2634;
   wire n_2635;
   wire n_2636;
   wire n_2637;
   wire n_2638;
   wire n_2639;
   wire n_2640;
   wire n_2641;
   wire n_2642;
   wire n_2643;
   wire n_2644;
   wire n_2645;
   wire n_2646;
   wire n_2647;
   wire n_2648;
   wire n_2649;
   wire n_2650;
   wire n_2651;
   wire n_2652;
   wire n_2653;
   wire n_2654;
   wire n_2655;
   wire n_2656;
   wire n_2657;
   wire n_2658;
   wire n_2659;
   wire n_2660;
   wire n_2661;
   wire n_2662;
   wire n_2663;
   wire n_2664;
   wire n_2665;
   wire n_2666;
   wire n_2667;
   wire n_2668;
   wire n_2669;
   wire n_2670;
   wire n_2671;
   wire n_2672;
   wire n_2673;
   wire n_2674;
   wire n_2675;
   wire n_2676;
   wire n_2677;
   wire n_2678;
   wire n_2679;
   wire n_2680;
   wire n_2681;
   wire n_2682;
   wire n_2683;
   wire n_2684;
   wire n_2685;
   wire n_2686;
   wire n_2687;
   wire n_2688;
   wire n_2689;
   wire n_2690;
   wire n_2691;
   wire n_2692;
   wire n_2693;
   wire n_2694;
   wire n_2695;
   wire n_2696;
   wire n_2697;
   wire n_2698;
   wire n_2699;
   wire n_2701;
   wire n_2702;
   wire n_2703;
   wire n_2704;
   wire n_2706;
   wire n_2708;
   wire n_2831;
   wire n_2834;
   wire n_2835;
   wire n_2836;

   INV_X1_50_SVT FE_PDC291_FE_OFN34_n_1383 (.A(FE_OFN34_n_1383),
	.Q(FE_PDN1444_FE_OFN34_n_1383));
   INV_X2_50_SVT FE_PDC290_FE_OFN34_n_1383 (.A(FE_PDN1444_FE_OFN34_n_1383),
	.Q(FE_PDN1443_FE_OFN34_n_1383));
   ANTENNA_50_SVT DIODE_9 (.I(DMEMRD[1]));
   ANTENNA_50_SVT DIODE_8 (.I(DMEMRD[5]));
   ANTENNA_50_SVT DIODE_7 (.I(DMEMRD[4]));
   ANTENNA_50_SVT DIODE_6 (.I(DMEMRD[7]));
   ANTENNA_50_SVT DIODE_5 (.I(DMEMRD[6]));
   ANTENNA_50_SVT DIODE_4 (.I(DMEMRD[2]));
   ANTENNA_50_SVT DIODE_3 (.I(DMEMRD[11]));
   ANTENNA_50_SVT DIODE_2 (.I(DMEMRD[22]));
   ANTENNA_50_SVT DIODE_1 (.I(DMEMRD[21]));
   CLKBUF_X2_50_SVT FE_OFC289_n_111 (.A(n_111),
	.Q(FE_OFN1442_n_111));
   CLKBUF_X2_50_SVT FE_OFC288_n_2619 (.A(n_2619),
	.Q(FE_OFN1441_n_2619));
   BUF_X2_50_SVT FE_OFC287_n_1389 (.A(n_1389),
	.Q(FE_OFN38_n_1389));
   INV_X2_50_SVT FE_OFC286_n_1427 (.A(n_1427),
	.Q(n_1426));
   BUF_X4_50_SVT FE_OFC285_n_1398 (.A(n_1398),
	.Q(FE_OFN46_n_1398));
   BUF_X4_50_SVT FE_OFC284_n_1392 (.A(n_1392),
	.Q(FE_OFN41_n_1392));
   BUF_X4_50_SVT FE_OFC283_n_1390 (.A(n_1390),
	.Q(FE_OFN39_n_1390));
   BUF_X4_50_SVT FE_OFC282_n_1396 (.A(n_1396),
	.Q(FE_OFN44_n_1396));
   BUF_X4_50_SVT FE_OFC281_n_1381 (.A(n_1381),
	.Q(FE_OFN33_n_1381));
   BUF_X4_50_SVT FE_OFC280_n_1422 (.A(n_1422),
	.Q(FE_OFN58_n_1422));
   BUF_X4_50_SVT FE_OFC279_n_1423 (.A(n_1423),
	.Q(FE_OFN59_n_1423));
   BUF_X4_50_SVT FE_OFC278_n_1393 (.A(n_1393),
	.Q(FE_OFN42_n_1393));
   BUF_X4_50_SVT FE_OFC277_n_1391 (.A(n_1391),
	.Q(FE_OFN40_n_1391));
   INVP2_X1_50_SVT FE_OFC276_n_1408 (.A(FE_OFN52_n_1408),
	.Q(n_1407));
   INV_X1_50_SVT FE_OFC275_n_1383 (.A(FE_PDN1443_FE_OFN34_n_1383),
	.Q(n_1382));
   INV_X1_50_SVT FE_OFC274_n_1395 (.A(FE_OFN43_n_1395),
	.Q(n_1394));
   INV_X1_50_SVT FE_OFC273_n_1331 (.A(FE_OFN25_n_1331),
	.Q(n_1388));
   INV_X1_50_SVT FE_OFC272_n_1419 (.A(FE_OFN57_n_1419),
	.Q(n_1418));
   CLKBUF_X6_50_SVT FE_OFC271_n_91 (.A(n_91),
	.Q(FE_OFN23_n_91));
   CLKBUF_X6_50_SVT FE_OFC270_n_76 (.A(n_76),
	.Q(FE_OFN77_n_76));
   CLKBUF_X6_50_SVT FE_OFC269_n_79 (.A(n_79),
	.Q(FE_OFN78_n_79));
   BUF_X4_50_SVT FE_OFC268_n_62 (.A(n_62),
	.Q(FE_OFN2_n_62));
   INV_X1_50_SVT FE_OFC267_DPATH_n_2548 (.A(DPATH_n_2548),
	.Q(n_2675));
   INV_X1_50_SVT FE_OFC266_DPATH_n_2538 (.A(DPATH_n_2538),
	.Q(n_2674));
   INV_X2_50_SVT FE_OFC265_n_132 (.A(FE_OFN103_n_132),
	.Q(n_131));
   INV_X2_50_SVT FE_OFC264_n_148 (.A(FE_OFN113_n_148),
	.Q(n_147));
   INV_X2_50_SVT FE_OFC263_n_115 (.A(FE_OFN92_n_115),
	.Q(n_114));
   INV_X2_50_SVT FE_OFC262_n_109 (.A(FE_OFN89_n_109),
	.Q(n_108));
   INV_X2_50_SVT FE_OFC261_n_103 (.A(FE_OFN86_n_103),
	.Q(n_102));
   INV_X2_50_SVT FE_OFC260_n_101 (.A(FE_OFN85_n_101),
	.Q(n_100));
   INV_X2_50_SVT FE_OFC259_OFN119_n_95 (.A(FE_OFN119_n_95),
	.Q(n_94));
   CLKBUF_X6_50_SVT CTS_cpc_drv_buf_00071 (.A(CTS_24),
	.Q(CTS_61));
   CLKBUF_X6_50_SVT CTS_cpc_drv_buf_00070 (.A(CTS_24),
	.Q(CTS_60));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00051 (.A(CTS_7),
	.Q(CTS_6));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00030 (.A(CTS_7),
	.Q(CTS_5));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00029 (.A(CTS_7),
	.Q(CTS_4));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00028 (.A(CTS_7),
	.Q(CTS_3));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00024 (.A(CTS_7),
	.Q(CTS_2));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00015 (.A(CTS_7),
	.Q(CTS_1));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00005 (.A(CTS_7),
	.Q(CTS_9));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00003 (.A(CTS_7),
	.Q(CTS_59));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00059 (.A(CLK),
	.Q(CTS_7));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00050 (.A(CTS_58),
	.Q(CTS_57));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00049 (.A(CTS_58),
	.Q(CTS_56));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00045 (.A(CTS_58),
	.Q(CTS_55));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00044 (.A(CTS_58),
	.Q(CTS_54));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00040 (.A(CTS_58),
	.Q(CTS_53));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00013 (.A(CTS_58),
	.Q(CTS_52));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00002 (.A(CTS_58),
	.Q(CTS_51));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00058 (.A(CLK),
	.Q(CTS_58));
   CLKBUF_X2_50_SVT CTS_ccl_a_buf_00048 (.A(CTS_25),
	.Q(CTS_24));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00047 (.A(CTS_25),
	.Q(CTS_23));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00046 (.A(CTS_25),
	.Q(CTS_27));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00037 (.A(CTS_25),
	.Q(CTS_50));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00057 (.A(CLK),
	.Q(CTS_25));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00043 (.A(CTS_49),
	.Q(CTS_48));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00042 (.A(CTS_49),
	.Q(CTS_47));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00041 (.A(CTS_49),
	.Q(CTS_46));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00036 (.A(CTS_49),
	.Q(CTS_45));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00021 (.A(CTS_49),
	.Q(CTS_44));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00008 (.A(CTS_49),
	.Q(CTS_43));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00007 (.A(CTS_49),
	.Q(CTS_42));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00056 (.A(CLK),
	.Q(CTS_49));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00039 (.A(CTS_20),
	.Q(CTS_19));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00038 (.A(CTS_20),
	.Q(CTS_18));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00032 (.A(CTS_20),
	.Q(CTS_17));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00018 (.A(CTS_20),
	.Q(CTS_16));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00017 (.A(CTS_20),
	.Q(CTS_15));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00016 (.A(CTS_20),
	.Q(CTS_22));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00014 (.A(CTS_20),
	.Q(CTS_41));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00055 (.A(CLK),
	.Q(CTS_20));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00035 (.A(CTS_12),
	.Q(CTS_11));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00027 (.A(CTS_12),
	.Q(CTS_10));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00026 (.A(CTS_12),
	.Q(CTS_14));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00012 (.A(CTS_12),
	.Q(CTS_40));
   CLKBUF_X2_50_SVT CTS_ccl_a_buf_00054 (.A(CLK),
	.Q(CTS_12));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00034 (.A(CTS_39),
	.Q(CTS_38));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00033 (.A(CTS_39),
	.Q(CTS_37));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00031 (.A(CTS_39),
	.Q(CTS_36));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00025 (.A(CTS_39),
	.Q(CTS_35));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00023 (.A(CTS_39),
	.Q(CTS_34));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00020 (.A(CTS_39),
	.Q(CTS_33));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00001 (.A(CTS_39),
	.Q(CTS_32));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00053 (.A(CLK),
	.Q(CTS_39));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00022 (.A(CTS_31),
	.Q(CTS_30));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00019 (.A(CTS_31),
	.Q(CTS_29));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00011 (.A(CTS_31),
	.Q(CTS_28));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00010 (.A(CTS_31),
	.Q(CTS_26));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00009 (.A(CTS_31),
	.Q(CTS_21));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00006 (.A(CTS_31),
	.Q(CTS_13));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00004 (.A(CTS_31),
	.Q(CTS_8));
   CLKBUF_X6_50_SVT CTS_ccl_a_buf_00052 (.A(CLK),
	.Q(CTS_31));
   INV_X1_50_SVT FE_OFC257_n_1348 (.A(n_1348),
	.Q(n_1347));
   INV_X1_50_SVT FE_OFC256_n_1335 (.A(n_1335),
	.Q(n_1334));
   INV_X1_50_SVT FE_OFC255_n_1350 (.A(n_1350),
	.Q(n_1349));
   INVP2_X1_50_SVT FE_OFC254_n_1338 (.A(n_1338),
	.Q(n_1337));
   CLKBUF_X4_50_SVT FE_OFC253_n_1380 (.A(n_1380),
	.Q(FE_OFN32_n_1380));
   CLKBUF_X4_50_SVT FE_OFC252_n_1442 (.A(n_1442),
	.Q(FE_OFN68_n_1442));
   CLKBUF_X4_50_SVT FE_OFC251_n_1441 (.A(n_1441),
	.Q(FE_OFN67_n_1441));
   INVP2_X1_50_SVT FE_OFC250_n_1438 (.A(FE_OFN65_n_1438),
	.Q(n_1437));
   CLKBUF_X4_50_SVT FE_OFC249_n_1438 (.A(n_1438),
	.Q(FE_OFN65_n_1438));
   CLKBUF_X4_50_SVT FE_OFC247_n_1379 (.A(n_1379),
	.Q(FE_OFN31_n_1379));
   INV_X4_50_SVT FE_OFC246_n_1332 (.A(n_1332),
	.Q(n_1372));
   CLKBUF_X4_50_SVT FE_OFC245_n_1377 (.A(n_1377),
	.Q(FE_OFN29_n_1377));
   CLKBUF_X4_50_SVT FE_OFC243_n_1408 (.A(n_1408),
	.Q(FE_OFN52_n_1408));
   INV_X1_50_SVT FE_OFC242_n_1436 (.A(FE_OFN64_n_1436),
	.Q(n_1435));
   BUF_X3_50_SVT FE_OFC241_n_1436 (.A(n_1436),
	.Q(FE_OFN64_n_1436));
   BUF_X3_50_SVT FE_OFC240_n_1371 (.A(n_1371),
	.Q(FE_OFN26_n_1371));
   INV_X1_50_SVT FE_OFC239_n_1440 (.A(n_1440),
	.Q(n_1439));
   BUF_X3_50_SVT FE_OFC238_n_1440 (.A(n_1440),
	.Q(FE_OFN66_n_1440));
   BUF_X3_50_SVT FE_OFC237_n_1386 (.A(n_1386),
	.Q(FE_OFN36_n_1386));
   INV_X2_50_SVT FE_OFC236_n_1403 (.A(n_1403),
	.Q(n_1402));
   CLKBUF_X4_50_SVT FE_OFC235_n_1409 (.A(n_1409),
	.Q(FE_OFN53_n_1409));
   CLKBUF_X4_50_SVT FE_OFC234_n_1413 (.A(n_1413),
	.Q(FE_OFN55_n_1413));
   CLKBUF_X4_50_SVT FE_OFC233_n_1411 (.A(n_1411),
	.Q(FE_OFN54_n_1411));
   CLKINV_X4_50_SVT FE_OFC231_n_1419 (.A(n_1419),
	.Q(FE_OFN57_n_1419));
   CLKBUF_X4_50_SVT FE_OFC230_n_1397 (.A(n_1397),
	.Q(FE_OFN45_n_1397));
   INV_X1_50_SVT FE_OFC229_n_1157 (.A(n_1157),
	.Q(n_1156));
   CLKBUF_X4_50_SVT FE_OFC221_n_1383 (.A(n_1383),
	.Q(FE_OFN34_n_1383));
   CLKINV_X4_50_SVT FE_OFC217_n_1415 (.A(FE_OFN56_n_1415),
	.Q(n_1414));
   INV_X1_50_SVT FE_OFC216_n_1415 (.A(n_1415),
	.Q(FE_OFN56_n_1415));
   CLKBUF_X4_50_SVT FE_OFC214_n_1395 (.A(n_1395),
	.Q(FE_OFN43_n_1395));
   INV_X2_50_SVT FE_OFC211_n_1425 (.A(FE_OFN60_n_1425),
	.Q(n_1424));
   INV_X1_50_SVT FE_OFC210_n_1425 (.A(n_1425),
	.Q(FE_OFN60_n_1425));
   INV_X2_50_SVT FE_OFC209_n_1432 (.A(FE_OFN63_n_1432),
	.Q(n_1431));
   INV_X2_50_SVT FE_OFC206_n_1376 (.A(FE_OFN28_n_1376),
	.Q(n_1375));
   INV_X2_50_SVT FE_OFC205_n_1374 (.A(FE_OFN27_n_1374),
	.Q(n_1373));
   INV_X2_50_SVT FE_OFC202_n_1429 (.A(FE_OFN62_n_1429),
	.Q(n_1428));
   INV_X1_50_SVT FE_OFC201_n_1385 (.A(FE_OFN35_n_1385),
	.Q(n_1384));
   CLKINV_X4_50_SVT FE_OFC193_n_1162 (.A(FE_OFN24_n_1162),
	.Q(n_1161));
   INV_X1_50_SVT FE_OFC192_n_28 (.A(n_28),
	.Q(n_27));
   INV_X2_50_SVT FE_OFC191_n_26 (.A(n_26),
	.Q(n_25));
   INVP2_X1_50_SVT FE_OFC190_n_24 (.A(n_24),
	.Q(n_23));
   CLKBUF_X6_50_SVT FE_OFC189_n_77 (.A(n_77),
	.Q(FE_OFN10_n_77));
   CLKBUF_X6_50_SVT FE_OFC188_n_89 (.A(n_89),
	.Q(FE_OFN21_n_89));
   CLKBUF_X6_50_SVT FE_OFC187_n_74 (.A(n_74),
	.Q(FE_OFN9_n_74));
   CLKBUF_X6_50_SVT FE_OFC186_n_84 (.A(n_84),
	.Q(FE_OFN16_n_84));
   CLKBUF_X6_50_SVT FE_OFC185_n_80 (.A(n_80),
	.Q(FE_OFN13_n_80));
   CLKBUF_X6_50_SVT FE_OFC184_n_90 (.A(n_90),
	.Q(FE_OFN22_n_90));
   CLKINV_X4_50_SVT FE_OFC183_n_1148 (.A(n_1148),
	.Q(n_1165));
   BUF_X6_50_SVT FE_OFC182_n_78 (.A(n_78),
	.Q(FE_OFN12_n_78));
   CLKBUF_X2_50_SVT FE_OFC181_n_82 (.A(n_82),
	.Q(FE_OFN79_n_82));
   CLKBUF_X4_50_SVT FE_OFC180_n_85 (.A(n_85),
	.Q(FE_OFN80_n_85));
   CLKBUF_X6_50_SVT FE_OFC179_n_67 (.A(n_67),
	.Q(FE_OFN4_n_67));
   CLKBUF_X6_50_SVT FE_OFC178_n_86 (.A(n_86),
	.Q(FE_OFN81_n_86));
   INV_X1_50_SVT FE_OFC173_DPATH_n_2496 (.A(DPATH_n_2496),
	.Q(n_2684));
   INV_X1_50_SVT FE_OFC172_DPATH_n_2498 (.A(DPATH_n_2498),
	.Q(n_2677));
   INV_X1_50_SVT FE_OFC171_DPATH_n_2508 (.A(DPATH_n_2508),
	.Q(n_2692));
   INV_X1_50_SVT FE_OFC170_DPATH_n_2550 (.A(DPATH_n_2550),
	.Q(n_2698));
   INV_X1_50_SVT FE_OFC169_DPATH_n_2552 (.A(DPATH_n_2552),
	.Q(n_2693));
   INV_X1_50_SVT FE_OFC168_DPATH_n_2512 (.A(DPATH_n_2512),
	.Q(n_2690));
   INV_X1_50_SVT FE_OFC167_DPATH_n_2514 (.A(DPATH_n_2514),
	.Q(n_2685));
   INV_X1_50_SVT FE_OFC166_DPATH_n_2544 (.A(DPATH_n_2544),
	.Q(n_2699));
   INV_X1_50_SVT FE_OFC165_DPATH_n_2530 (.A(DPATH_n_2530),
	.Q(n_2681));
   INV_X1_50_SVT FE_OFC164_DPATH_n_2542 (.A(DPATH_n_2542),
	.Q(n_2689));
   INV_X1_50_SVT FE_OFC163_DPATH_n_2534 (.A(DPATH_n_2534),
	.Q(n_2678));
   INV_X1_50_SVT FE_OFC162_DPATH_n_2506 (.A(DPATH_n_2506),
	.Q(n_2701));
   INV_X1_50_SVT FE_OFC161_DPATH_n_2502 (.A(DPATH_n_2502),
	.Q(n_2694));
   INV_X1_50_SVT FE_OFC160_DPATH_B_31 (.A(DPATH_B_31_),
	.Q(n_1149));
   INV_X1_50_SVT FE_OFC159_DPATH_n_2556 (.A(DPATH_n_2556),
	.Q(n_2702));
   INV_X1_50_SVT FE_OFC158_DPATH_n_2554 (.A(DPATH_n_2554),
	.Q(n_2687));
   INV_X1_50_SVT FE_OFC157_DPATH_n_2536 (.A(DPATH_n_2536),
	.Q(n_2676));
   INV_X1_50_SVT FE_OFC156_DPATH_n_2520 (.A(DPATH_n_2520),
	.Q(n_2696));
   INV_X1_50_SVT FE_OFC155_DPATH_n_2532 (.A(DPATH_n_2532),
	.Q(n_2680));
   INV_X1_50_SVT FE_OFC154_DPATH_n_2540 (.A(DPATH_n_2540),
	.Q(n_2688));
   INV_X1_50_SVT FE_OFC153_DPATH_n_2546 (.A(DPATH_n_2546),
	.Q(n_2679));
   INV_X1_50_SVT FE_OFC152_DPATH_n_2516 (.A(DPATH_n_2516),
	.Q(n_2682));
   INV_X1_50_SVT FE_OFC151_DPATH_n_2526 (.A(DPATH_n_2526),
	.Q(n_2673));
   INV_X1_50_SVT FE_OFC150_DPATH_n_2522 (.A(DPATH_n_2522),
	.Q(n_2695));
   INV_X1_50_SVT FE_OFC149_DPATH_n_2504 (.A(DPATH_n_2504),
	.Q(n_2683));
   INV_X1_50_SVT FE_OFC148_DPATH_n_2528 (.A(DPATH_n_2528),
	.Q(n_2686));
   INV_X1_50_SVT FE_OFC147_DPATH_n_2524 (.A(DPATH_n_2524),
	.Q(n_2691));
   INV_X1_50_SVT FE_OFC146_DPATH_n_2510 (.A(DPATH_n_2510),
	.Q(n_2703));
   INV_X1_50_SVT FE_OFC145_DPATH_n_2518 (.A(DPATH_n_2518),
	.Q(n_2704));
   INV_X1_50_SVT FE_OFC142_DPATH_n_2500 (.A(DPATH_n_2500),
	.Q(n_2697));
   INV_X2_50_SVT FE_OFC141_n_140 (.A(FE_OFN108_n_140),
	.Q(n_139));
   CLKBUF_X2_50_SVT FE_OFC140_n_140 (.A(n_140),
	.Q(FE_OFN108_n_140));
   CLKBUF_X2_50_SVT FE_OFC139_n_128 (.A(n_128),
	.Q(FE_OFN101_n_128));
   INV_X2_50_SVT FE_OFC138_n_93 (.A(FE_OFN82_n_93),
	.Q(n_92));
   CLKBUF_X2_50_SVT FE_OFC136_n_132 (.A(n_132),
	.Q(FE_OFN103_n_132));
   CLKBUF_X4_50_SVT FE_OFC134_n_148 (.A(n_148),
	.Q(FE_OFN113_n_148));
   CLKBUF_X4_50_SVT FE_OFC131_n_115 (.A(n_115),
	.Q(FE_OFN92_n_115));
   INV_X2_50_SVT FE_OFC129_n_113 (.A(FE_OFN91_n_113),
	.Q(n_112));
   CLKBUF_X2_50_SVT FE_OFC128_n_113 (.A(n_113),
	.Q(FE_OFN91_n_113));
   CLKBUF_X4_50_SVT FE_OFC126_n_109 (.A(n_109),
	.Q(FE_OFN89_n_109));
   CLKBUF_X2_50_SVT FE_OFC124_n_103 (.A(n_103),
	.Q(FE_OFN86_n_103));
   CLKBUF_X2_50_SVT FE_OFC122_n_101 (.A(n_101),
	.Q(FE_OFN85_n_101));
   CLKBUF_X2_50_SVT FE_OFC120_95 (.A(n_95),
	.Q(FE_OFN119_n_95));
   CLKBUF_X2_50_SVT FE_OFC118_n_1198 (.A(n_1198),
	.Q(FE_OFN118_n_1198));
   CLKBUF_X2_50_SVT FE_OFC117_n_154 (.A(n_154),
	.Q(FE_OFN117_n_154));
   INV_X2_50_SVT FE_OFC116_n_152 (.A(FE_OFN115_n_152),
	.Q(FE_OFN116_n_152));
   INV_X1_50_SVT FE_OFC115_n_152 (.A(n_152),
	.Q(FE_OFN115_n_152));
   CLKBUF_X2_50_SVT FE_OFC114_n_150 (.A(n_150),
	.Q(FE_OFN114_n_150));
   CLKBUF_X2_50_SVT FE_OFC112_n_146 (.A(n_146),
	.Q(FE_OFN112_n_146));
   CLKBUF_X2_50_SVT FE_OFC111_n_144 (.A(n_144),
	.Q(FE_OFN111_n_144));
   INV_X2_50_SVT FE_OFC110_n_142 (.A(FE_OFN109_n_142),
	.Q(FE_OFN110_n_142));
   INV_X1_50_SVT FE_OFC109_n_142 (.A(n_142),
	.Q(FE_OFN109_n_142));
   CLKBUF_X2_50_SVT FE_OFC107_n_138 (.A(n_138),
	.Q(FE_OFN107_n_138));
   CLKBUF_X2_50_SVT FE_OFC106_n_136 (.A(n_136),
	.Q(FE_OFN106_n_136));
   INV_X2_50_SVT FE_OFC105_n_134 (.A(FE_OFN104_n_134),
	.Q(FE_OFN105_n_134));
   INV_X1_50_SVT FE_OFC104_n_134 (.A(n_134),
	.Q(FE_OFN104_n_134));
   CLKBUF_X2_50_SVT FE_OFC102_n_130 (.A(n_130),
	.Q(FE_OFN102_n_130));
   CLKBUF_X2_50_SVT FE_OFC100_n_127 (.A(n_127),
	.Q(FE_OFN100_n_127));
   INV_X2_50_SVT FE_OFC99_n_125 (.A(FE_OFN98_n_125),
	.Q(FE_OFN99_n_125));
   INV_X1_50_SVT FE_OFC98_n_125 (.A(n_125),
	.Q(FE_OFN98_n_125));
   CLKBUF_X2_50_SVT FE_OFC97_n_123 (.A(n_123),
	.Q(FE_OFN97_n_123));
   CLKBUF_X2_50_SVT FE_OFC96_n_121 (.A(n_121),
	.Q(FE_OFN96_n_121));
   INV_X2_50_SVT FE_OFC95_n_119 (.A(FE_OFN94_n_119),
	.Q(FE_OFN95_n_119));
   INV_X1_50_SVT FE_OFC94_n_119 (.A(n_119),
	.Q(FE_OFN94_n_119));
   CLKBUF_X2_50_SVT FE_OFC93_n_117 (.A(n_117),
	.Q(FE_OFN93_n_117));
   CLKBUF_X2_50_SVT FE_OFC90_n_111 (.A(FE_OFN1442_n_111),
	.Q(FE_OFN90_n_111));
   CLKBUF_X2_50_SVT FE_OFC88_n_107 (.A(n_107),
	.Q(FE_OFN88_n_107));
   CLKBUF_X2_50_SVT FE_OFC87_n_105 (.A(n_105),
	.Q(FE_OFN87_n_105));
   CLKBUF_X2_50_SVT FE_OFC84_n_99 (.A(n_99),
	.Q(FE_OFN84_n_99));
   CLKBUF_X2_50_SVT FE_OFC83_n_97 (.A(n_97),
	.Q(FE_OFN83_n_97));
   CLKBUF_X2_50_SVT FE_OFC82_n_93 (.A(n_93),
	.Q(FE_OFN82_n_93));
   BUF_X6_50_SVT FE_OFC76_n_75 (.A(n_75),
	.Q(FE_OFN76_n_75));
   BUF_X6_50_SVT FE_OFC75_n_73 (.A(n_73),
	.Q(FE_OFN75_n_73));
   CLKBUF_X2_50_SVT FE_OFC74_n_72 (.A(n_72),
	.Q(FE_OFN74_n_72));
   BUF_X4_50_SVT FE_OFC73_n_1449 (.A(n_1449),
	.Q(FE_OFN73_n_1449));
   BUF_X4_50_SVT FE_OFC72_n_1448 (.A(n_1448),
	.Q(FE_OFN72_n_1448));
   BUF_X4_50_SVT FE_OFC69_n_1443 (.A(n_1443),
	.Q(FE_OFN69_n_1443));
   CLKBUF_X4_50_SVT FE_OFC63_n_1432 (.A(n_1432),
	.Q(FE_OFN63_n_1432));
   CLKBUF_X6_50_SVT FE_OFC62_n_1429 (.A(n_1429),
	.Q(FE_OFN62_n_1429));
   BUF_X4_50_SVT FE_OFC49_n_1404 (.A(n_1404),
	.Q(FE_OFN49_n_1404));
   CLKBUF_X6_50_SVT FE_OFC48_n_1401 (.A(n_1401),
	.Q(FE_OFN48_n_1401));
   BUF_X4_50_SVT FE_OFC47_n_1400 (.A(n_1400),
	.Q(FE_OFN47_n_1400));
   CLKBUF_X4_50_SVT FE_OFC35_n_1385 (.A(n_1385),
	.Q(FE_OFN35_n_1385));
   CLKBUF_X4_50_SVT FE_OFC28_n_1376 (.A(n_1376),
	.Q(FE_OFN28_n_1376));
   CLKBUF_X4_50_SVT FE_OFC27_n_1374 (.A(n_1374),
	.Q(FE_OFN27_n_1374));
   CLKBUF_X4_50_SVT FE_OFC25_n_1331 (.A(n_1331),
	.Q(FE_OFN25_n_1331));
   CLKBUF_X2_50_SVT FE_OFC24_n_1162 (.A(n_1162),
	.Q(FE_OFN24_n_1162));
   CLKBUF_X6_50_SVT FE_OFC19_n_88 (.A(n_88),
	.Q(FE_OFN19_n_88));
   CLKBUF_X6_50_SVT FE_OFC17_n_87 (.A(n_87),
	.Q(FE_OFN17_n_87));
   BUF_X6_50_SVT FE_OFC15_n_83 (.A(n_83),
	.Q(FE_OFN15_n_83));
   BUF_X6_50_SVT FE_OFC8_n_71 (.A(n_71),
	.Q(FE_OFN8_n_71));
   CLKBUF_X6_50_SVT FE_OFC6_n_70 (.A(n_70),
	.Q(FE_OFN6_n_70));
   BUF_X6_50_SVT FE_OFC5_n_69 (.A(n_69),
	.Q(FE_OFN5_n_69));
   BUF_X6_50_SVT FE_OFC3_n_64 (.A(n_64),
	.Q(FE_OFN3_n_64));
   BUF_X6_50_SVT FE_OFC0_n_2 (.A(n_2),
	.Q(FE_OFN0_n_2));
   INV_X4_50_SVT g24167 (.A(RST),
	.Q(n_2672));
   NAND2_A_NAND2_X0_50_SVT g78452__2398 (.A0N(WRDATA[15]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2526));
   NAND2_A_NAND2_X0_50_SVT g78453__5107 (.A0N(WRDATA[12]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2532));
   MUX2_X0_50_SVT g78454__6260 (.A(INSTR[30]),
	.B(WRDATA[10]),
	.Q(DPATH_n_2536),
	.S0(n_1356));
   MUX2_X0_50_SVT g78455__4319 (.A(n_2831),
	.B(WRDATA[0]),
	.Q(DPATH_n_2556),
	.S0(n_1356));
   NAND2_A_NAND2_X0_50_SVT g78456__8428 (.A0N(WRDATA[28]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2500));
   NAND2_A_NAND2_X0_50_SVT g78457__5526 (.A0N(WRDATA[27]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2502));
   NAND4_X2_50_SVT g78458__6783 (.A(n_2669),
	.B(n_2228),
	.C(n_1626),
	.D(n_1621),
	.Q(WRDATA[12]));
   NAND4_X2_50_SVT g78459__3680 (.A(n_2668),
	.B(n_2221),
	.C(n_1512),
	.D(n_1503),
	.Q(WRDATA[10]));
   NAND4_X2_50_SVT g78460__1617 (.A(n_2670),
	.B(n_2237),
	.C(n_1791),
	.D(n_1795),
	.Q(WRDATA[15]));
   NAND4_X2_50_SVT g78461__2802 (.A(n_2671),
	.B(n_2238),
	.C(n_1831),
	.D(n_1830),
	.Q(WRDATA[0]));
   MUX2_X0_50_SVT g78462__1705 (.A(DPATH_n_5229),
	.B(WRDATA[1]),
	.Q(DPATH_n_2554),
	.S0(n_1356));
   NAND2_A_NAND2_X0_50_SVT g78463__5122 (.A0N(WRDATA[16]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2524));
   NAND2_A_NAND2_X0_50_SVT g78464__8246 (.A0N(WRDATA[14]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2528));
   NAND2_A_NAND2_X0_50_SVT g78465__7098 (.A0N(WRDATA[11]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2534));
   MUX2_X0_50_SVT g78466__6131 (.A(INSTR[29]),
	.B(WRDATA[9]),
	.Q(DPATH_n_2538),
	.S0(n_1356));
   MUX2_X0_50_SVT g78467__1881 (.A(INSTR[28]),
	.B(WRDATA[8]),
	.Q(DPATH_n_2540),
	.S0(n_1356));
   NAND2_A_NAND2_X0_50_SVT g78468__5115 (.A0N(WRDATA[26]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2504));
   NAND2_A_NAND2_X0_50_SVT g78469__7482 (.A0N(WRDATA[18]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2520));
   NAND2_A_NAND2_X0_50_SVT g78470__4733 (.A0N(WRDATA[23]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2510));
   NAND2_A_NAND2_X0_50_SVT g78471__6161 (.A0N(WRDATA[21]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2514));
   NAND2_A_NAND2_X0_50_SVT g78472__9315 (.A0N(WRDATA[29]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2498));
   NAND2_A_NAND2_X0_50_SVT g78473__9945 (.A0N(WRDATA[22]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2512));
   NAND2_A_NAND2_X0_50_SVT g78474__2883 (.A0N(WRDATA[24]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2508));
   NAND2_A_NAND2_X0_50_SVT g78475__2346 (.A0N(WRDATA[30]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2496));
   NAND2_A_NAND2_X0_50_SVT g78476__1666 (.A0N(WRDATA[20]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2516));
   NAND2_A_NAND2_X0_50_SVT g78477__7410 (.A0N(WRDATA[25]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2506));
   NAND2_A_NAND2_X0_50_SVT g78478__6417 (.A0N(WRDATA[17]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2522));
   NAND2_A_NAND2_X0_50_SVT g78479__5477 (.A0N(WRDATA[19]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2518));
   NAND2_A_NAND2_X0_50_SVT g78480__2398 (.A0N(WRDATA[13]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_n_2530));
   NAND2_A_NAND2_X0_50_SVT g78481__5107 (.A0N(WRDATA[31]),
	.A1N(n_1356),
	.B0(n_1330),
	.Q(DPATH_B_31_));
   MUX2_X0_50_SVT g78482__6260 (.A(INSTR[27]),
	.B(WRDATA[7]),
	.Q(DPATH_n_2542),
	.S0(n_1356));
   MUX2_X0_50_SVT g78483__4319 (.A(INSTR[26]),
	.B(WRDATA[6]),
	.Q(DPATH_n_2544),
	.S0(n_1356));
   MUX2_X0_50_SVT g78484__8428 (.A(INSTR[25]),
	.B(WRDATA[5]),
	.Q(DPATH_n_2546),
	.S0(n_1356));
   MUX2_X0_50_SVT g78485__5526 (.A(DPATH_n_5226),
	.B(WRDATA[4]),
	.Q(DPATH_n_2548),
	.S0(n_1356));
   MUX2_X0_50_SVT g78486__6783 (.A(DPATH_n_5227),
	.B(WRDATA[3]),
	.Q(DPATH_n_2550),
	.S0(n_1356));
   MUX2_X0_50_SVT g78487__3680 (.A(DPATH_n_5228),
	.B(WRDATA[2]),
	.Q(DPATH_n_2552),
	.S0(n_1356));
   NOR2_A_NAND3_X2_50_SVT g78488__1617 (.AN(n_2407),
	.BN(n_2659),
	.C(n_1854),
	.D(n_2483),
	.Q(WRDATA[1]));
   NOR2_A_NAND3_X1_50_SVT g78489__2802 (.AN(n_2466),
	.BN(n_2662),
	.C(n_2180),
	.D(n_2449),
	.Q(WRDATA[9]));
   NOR2_A_NAND3_X1_50_SVT g78490__1705 (.AN(n_2455),
	.BN(n_2667),
	.C(n_2127),
	.D(n_2485),
	.Q(WRDATA[8]));
   NOR2_A_NAND3_X2_50_SVT g78491__5122 (.AN(n_2396),
	.BN(n_2654),
	.C(n_1897),
	.D(n_2481),
	.Q(WRDATA[28]));
   NOR2_A_NAND3_X1_50_SVT g78492__8246 (.AN(n_2403),
	.BN(n_2658),
	.C(n_1842),
	.D(n_2482),
	.Q(WRDATA[16]));
   NOR2_A_NAND3_X1_50_SVT g78493__7098 (.AN(n_2400),
	.BN(n_2657),
	.C(n_1806),
	.D(n_2480),
	.Q(DPATH_A_31_));
   NOR2_A_NAND3_X1_50_SVT g78494__6131 (.AN(n_2381),
	.BN(n_2656),
	.C(n_1740),
	.D(n_2479),
	.Q(WRDATA[14]));
   NOR2_A_NAND3_X2_50_SVT g78495__1881 (.AN(n_2350),
	.BN(n_2655),
	.C(n_1696),
	.D(n_2478),
	.Q(WRDATA[27]));
   NOR2_A_NAND3_X1_50_SVT g78496__5115 (.AN(n_2348),
	.BN(n_2660),
	.C(n_1570),
	.D(n_2477),
	.Q(WRDATA[11]));
   NAND4_X2_50_SVT g78497__7482 (.A(n_2663),
	.B(n_2445),
	.C(n_2484),
	.D(n_2193),
	.Q(WRDATA[26]));
   INV_A_OAI211_X2_50_SVT g78498__4733 (.A0(n_1435),
	.A1N(DPATH_RF_MEMORY_21__12_),
	.B0(n_2647),
	.C0(n_2603),
	.Q(DPATH_n_2402));
   INV_A_OAI211_X2_50_SVT g78499__6161 (.A0(n_1439),
	.A1N(DPATH_RF_MEMORY_19__10_),
	.B0(n_2651),
	.C0(n_2574),
	.Q(DPATH_n_2404));
   INV_A_OAI211_X2_50_SVT g78500__9315 (.A0(n_1437),
	.A1N(DPATH_RF_MEMORY_22__28_),
	.B0(n_2648),
	.C0(n_2599),
	.Q(DPATH_n_2386));
   INV_A_OAI211_X2_50_SVT g78501__9945 (.A0(n_1407),
	.A1N(DPATH_RF_MEMORY_20__27_),
	.B0(n_2646),
	.C0(n_2598),
	.Q(DPATH_n_2387));
   INV_A_OAI211_X2_50_SVT g78502__2883 (.A0(n_1437),
	.A1N(DPATH_RF_MEMORY_22__20_),
	.B0(n_2645),
	.C0(n_2597),
	.Q(DPATH_n_2394));
   INV_A_OAI211_X2_50_SVT g78503__2346 (.A0(n_1407),
	.A1N(DPATH_RF_MEMORY_20__19_),
	.B0(n_2644),
	.C0(n_2596),
	.Q(DPATH_n_2395));
   AOI221_X1_50_SVT g78504__1666 (.A0(DPATH_RF_MEMORY_21__0_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__0_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2661),
	.Q(n_2671));
   AOI221_X1_50_SVT g78505__7410 (.A0(DPATH_RF_MEMORY_20__15_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__15_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2666),
	.Q(n_2670));
   AOI221_X1_50_SVT g78506__6417 (.A0(DPATH_RF_MEMORY_20__12_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__12_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2665),
	.Q(n_2669));
   AOI221_X1_50_SVT g78507__5477 (.A0(DPATH_RF_MEMORY_20__10_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__10_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2664),
	.Q(n_2668));
   NAND4_X2_50_SVT g78508__2398 (.A(n_2626),
	.B(n_2528),
	.C(n_2453),
	.D(n_2081),
	.Q(DPATH_n_2406));
   NAND4_X2_50_SVT g78509__5107 (.A(n_2625),
	.B(n_2526),
	.C(n_2486),
	.D(n_2063),
	.Q(DPATH_n_2407));
   NAND4_X2_50_SVT g78510__6260 (.A(n_2623),
	.B(n_2525),
	.C(n_2446),
	.D(n_2041),
	.Q(DPATH_n_2408));
   NAND4_X2_50_SVT g78511__4319 (.A(n_2621),
	.B(n_2522),
	.C(n_2436),
	.D(n_1986),
	.Q(DPATH_n_2411));
   NAND4_X2_50_SVT g78512__8428 (.A(FE_OFN1441_n_2619),
	.B(n_2521),
	.C(n_2427),
	.D(n_1940),
	.Q(DPATH_n_2414));
   NAND4_X2_50_SVT g78513__5526 (.A(n_2615),
	.B(n_2510),
	.C(n_2397),
	.D(n_1769),
	.Q(DPATH_n_2384));
   NAND4_X2_50_SVT g78514__6783 (.A(n_2614),
	.B(n_2507),
	.C(n_2391),
	.D(n_1750),
	.Q(DPATH_n_2385));
   INV_A_OAI211_X2_50_SVT g78515__3680 (.A0(n_1388),
	.A1N(DPATH_RF_MEMORY_22__4_),
	.B0(n_2649),
	.C0(n_2594),
	.Q(WRDATA[4]));
   INV_A_OAI211_X2_50_SVT g78516__1617 (.A0(FE_OFN60_n_1425),
	.A1N(DPATH_RF_MEMORY_21__31_),
	.B0(n_2650),
	.C0(n_2595),
	.Q(WRDATA[31]));
   NAND4_X2_50_SVT g78517__2802 (.A(n_2622),
	.B(n_2527),
	.C(n_2448),
	.D(n_2036),
	.Q(WRDATA[7]));
   NAND4_X2_50_SVT g78518__1705 (.A(n_2620),
	.B(n_2523),
	.C(n_2438),
	.D(n_1982),
	.Q(WRDATA[6]));
   NAND4_X2_50_SVT g78519__5122 (.A(n_2519),
	.B(n_2618),
	.C(n_2418),
	.D(n_1887),
	.Q(WRDATA[3]));
   NAND4_X2_50_SVT g78520__8246 (.A(n_2612),
	.B(n_2524),
	.C(n_2375),
	.D(n_1765),
	.Q(WRDATA[30]));
   NAND4_X2_50_SVT g78521__7098 (.A(n_2617),
	.B(n_2517),
	.C(n_2413),
	.D(n_1865),
	.Q(WRDATA[2]));
   NAND4_X2_50_SVT g78522__6131 (.A(n_2616),
	.B(n_2515),
	.C(n_2408),
	.D(n_1807),
	.Q(WRDATA[24]));
   INV_A_OAI211_X2_50_SVT g78523__1881 (.A0(n_1388),
	.A1N(DPATH_RF_MEMORY_22__20_),
	.B0(n_2652),
	.C0(n_2602),
	.Q(WRDATA[20]));
   INV_A_OAI211_X2_50_SVT g78524__5115 (.A0(n_1388),
	.A1N(DPATH_RF_MEMORY_22__23_),
	.B0(n_2653),
	.C0(n_2600),
	.Q(WRDATA[23]));
   NAND4_X2_50_SVT g78525__7482 (.A(n_2642),
	.B(n_2217),
	.C(n_2146),
	.D(n_1465),
	.Q(DPATH_n_2403));
   NAND4_X2_50_SVT g78526__4733 (.A(n_2610),
	.B(n_2499),
	.C(n_2369),
	.D(n_1636),
	.Q(DPATH_n_2391));
   NAND4_X2_50_SVT g78527__6161 (.A(n_2609),
	.B(n_2498),
	.C(n_2366),
	.D(n_1614),
	.Q(DPATH_n_2392));
   NAND4_X2_50_SVT g78528__9315 (.A(n_2608),
	.B(n_2497),
	.C(n_2363),
	.D(n_1597),
	.Q(DPATH_n_2393));
   NAND4_X2_50_SVT g78529__9945 (.A(n_2606),
	.B(n_2490),
	.C(n_2346),
	.D(n_1523),
	.Q(DPATH_n_2397));
   NAND4_X2_50_SVT g78530__2883 (.A(n_2605),
	.B(n_2489),
	.C(n_2343),
	.D(n_1502),
	.Q(DPATH_n_2398));
   NAND4_X2_50_SVT g78531__2346 (.A(n_2604),
	.B(n_2488),
	.C(n_2340),
	.D(n_1482),
	.Q(DPATH_n_2399));
   NAND4_X2_50_SVT g78532__1666 (.A(n_2627),
	.B(n_2530),
	.C(n_2475),
	.D(n_2191),
	.Q(DPATH_n_2400));
   NAND4_X2_50_SVT g78533__7410 (.A(n_2643),
	.B(n_2218),
	.C(n_2182),
	.D(n_1454),
	.Q(DPATH_n_2401));
   NAND4_X2_50_SVT g78534__6417 (.A(n_2613),
	.B(n_2503),
	.C(n_2380),
	.D(n_1693),
	.Q(DPATH_n_2388));
   NAND4_X2_50_SVT g78535__5477 (.A(n_2641),
	.B(n_2216),
	.C(n_2110),
	.D(n_1459),
	.Q(DPATH_n_2405));
   NAND4_X2_50_SVT g78536__2398 (.A(n_2640),
	.B(n_2215),
	.C(n_2054),
	.D(n_1464),
	.Q(DPATH_n_2409));
   NAND4_X2_50_SVT g78537__5107 (.A(n_2638),
	.B(n_2213),
	.C(n_2017),
	.D(n_1456),
	.Q(DPATH_n_2410));
   NAND4_X2_50_SVT g78538__6260 (.A(n_2637),
	.B(n_2212),
	.C(n_1978),
	.D(n_1466),
	.Q(DPATH_n_2412));
   NAND4_X2_50_SVT g78539__4319 (.A(n_2636),
	.B(n_2211),
	.C(n_1964),
	.D(n_1463),
	.Q(DPATH_n_2413));
   NAND4_X2_50_SVT g78540__8428 (.A(n_2631),
	.B(n_2206),
	.C(n_1684),
	.D(n_1455),
	.Q(DPATH_n_2389));
   NAND4_X2_50_SVT g78541__5526 (.A(n_2630),
	.B(n_2205),
	.C(n_1667),
	.D(n_1453),
	.Q(DPATH_n_2390));
   NAND4_X2_50_SVT g78542__6783 (.A(n_2629),
	.B(n_2204),
	.C(n_1554),
	.D(n_1457),
	.Q(DPATH_n_2396));
   NAND4_X2_50_SVT g78543__3680 (.A(n_2633),
	.B(n_2203),
	.C(n_1929),
	.D(n_1461),
	.Q(WRDATA[18]));
   NAND4_X2_50_SVT g78544__1617 (.A(n_2611),
	.B(n_2502),
	.C(n_2412),
	.D(n_1653),
	.Q(WRDATA[13]));
   NAND4_X2_50_SVT g78545__2802 (.A(n_2628),
	.B(n_2491),
	.C(n_2344),
	.D(n_2199),
	.Q(WRDATA[21]));
   NAND4_X2_50_SVT g78546__1705 (.A(n_2634),
	.B(n_2210),
	.C(n_1962),
	.D(n_1460),
	.Q(WRDATA[5]));
   NAND4_X2_50_SVT g78547__5122 (.A(n_2635),
	.B(n_2209),
	.C(n_1970),
	.D(n_1452),
	.Q(WRDATA[25]));
   NAND4_X2_50_SVT g78548__8246 (.A(n_2632),
	.B(n_2207),
	.C(n_1885),
	.D(n_1458),
	.Q(WRDATA[17]));
   NAND4_X2_50_SVT g78549__7098 (.A(n_2624),
	.B(n_2494),
	.C(n_2468),
	.D(n_2032),
	.Q(WRDATA[29]));
   NAND4_X2_50_SVT g78550__6131 (.A(n_2639),
	.B(n_2214),
	.C(n_2033),
	.D(n_1462),
	.Q(WRDATA[19]));
   NAND4_X2_50_SVT g78551__1881 (.A(n_2607),
	.B(n_2501),
	.C(n_2368),
	.D(n_1587),
	.Q(WRDATA[22]));
   INV_A_OAI211_X2_50_SVT g78552__5115 (.A0(n_1428),
	.A1N(DPATH_RF_MEMORY_15__8_),
	.B0(n_2591),
	.C0(n_2119),
	.Q(n_2667));
   NAND4_X2_50_SVT g78553__7482 (.A(n_2508),
	.B(n_2398),
	.C(n_1780),
	.D(n_1761),
	.Q(n_2666));
   NAND4_X2_50_SVT g78554__4733 (.A(n_2495),
	.B(n_2364),
	.C(n_1607),
	.D(n_1588),
	.Q(n_2665));
   NAND4_X2_50_SVT g78555__6161 (.A(n_2533),
	.B(n_2341),
	.C(n_1489),
	.D(n_1470),
	.Q(n_2664));
   AOI211_X2_50_SVT g78556__9315 (.A0(DPATH_RF_MEMORY_16__26_),
	.A1(FE_OFN43_n_1395),
	.B0(n_2170),
	.C0(n_2592),
	.Q(n_2663));
   INV_A_OAI211_X1_50_SVT g78557__9945 (.A0(n_1428),
	.A1N(DPATH_RF_MEMORY_15__9_),
	.B0(n_2593),
	.C0(n_2174),
	.Q(n_2662));
   NAND4_X2_50_SVT g78558__2883 (.A(n_2512),
	.B(n_2405),
	.C(n_1824),
	.D(n_1815),
	.Q(n_2661));
   INV_A_OAI211_X2_50_SVT g78559__2346 (.A0(n_1402),
	.A1N(DPATH_RF_MEMORY_7__11_),
	.B0(n_2584),
	.C0(n_1564),
	.Q(n_2660));
   INV_A_OAI211_X2_50_SVT g78560__1666 (.A0(n_1375),
	.A1N(DPATH_RF_MEMORY_1__1_),
	.B0(n_2589),
	.C0(n_1852),
	.Q(n_2659));
   INV_A_OAI211_X2_50_SVT g78561__7410 (.A0(n_1402),
	.A1N(DPATH_RF_MEMORY_7__16_),
	.B0(n_2588),
	.C0(n_2201),
	.Q(n_2658));
   INV_A_OAI211_X2_50_SVT g78562__6417 (.A0(n_1433),
	.A1N(DPATH_RF_MEMORY_2__31_),
	.B0(n_2587),
	.C0(n_1802),
	.Q(n_2657));
   INV_A_OAI211_X1_50_SVT g78563__5477 (.A0(n_1402),
	.A1N(DPATH_RF_MEMORY_7__14_),
	.B0(n_2586),
	.C0(n_1732),
	.Q(n_2656));
   INV_A_OAI211_X2_50_SVT g78564__2398 (.A0(n_1382),
	.A1N(DPATH_RF_MEMORY_9__27_),
	.B0(n_2585),
	.C0(n_1665),
	.Q(n_2655));
   INV_A_OAI211_X2_50_SVT g78565__5107 (.A0(n_1375),
	.A1N(DPATH_RF_MEMORY_1__28_),
	.B0(n_2590),
	.C0(n_1879),
	.Q(n_2654));
   AOI221_X1_50_SVT g78566__6260 (.A0(DPATH_RF_MEMORY_17__23_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__23_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2577),
	.Q(n_2653));
   AOI221_X1_50_SVT g78567__4319 (.A0(DPATH_RF_MEMORY_17__20_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__20_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2580),
	.Q(n_2652));
   AOI221_X1_50_SVT g78568__8428 (.A0(DPATH_RF_MEMORY_17__10_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__10_),
	.B1(n_1386),
	.C0(n_2581),
	.Q(n_2651));
   AOI221_X1_50_SVT g78569__5526 (.A0(DPATH_RF_MEMORY_18__31_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__31_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2583),
	.Q(n_2650));
   AOI221_X1_50_SVT g78570__6783 (.A0(DPATH_RF_MEMORY_17__4_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__4_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2579),
	.Q(n_2649));
   AOI221_X1_50_SVT g78571__3680 (.A0(DPATH_RF_MEMORY_17__28_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__28_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2578),
	.Q(n_2648));
   AOI221_X1_50_SVT g78572__1617 (.A0(DPATH_RF_MEMORY_17__12_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__12_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2582),
	.Q(n_2647));
   AOI221_X1_50_SVT g78573__2802 (.A0(DPATH_RF_MEMORY_17__27_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__27_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2576),
	.Q(n_2646));
   AOI221_X1_50_SVT g78574__1705 (.A0(DPATH_RF_MEMORY_17__20_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__20_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2575),
	.Q(n_2645));
   AOI221_X1_50_SVT g78575__5122 (.A0(DPATH_RF_MEMORY_17__19_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__19_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2601),
	.Q(n_2644));
   AOI211_X2_50_SVT g78576__8246 (.A0(DPATH_RF_MEMORY_18__13_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2474),
	.C0(n_2552),
	.Q(n_2643));
   AOI211_X2_50_SVT g78577__7098 (.A0(DPATH_RF_MEMORY_18__11_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2467),
	.C0(n_2572),
	.Q(n_2642));
   AOI211_X2_50_SVT g78578__6131 (.A0(DPATH_RF_MEMORY_18__9_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2458),
	.C0(n_2571),
	.Q(n_2641));
   AOI211_X2_50_SVT g78579__1881 (.A0(DPATH_RF_MEMORY_18__5_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2444),
	.C0(n_2570),
	.Q(n_2640));
   AOI211_X1_50_SVT g78580__5115 (.A0(DPATH_RF_MEMORY_18__19_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2442),
	.C0(n_2568),
	.Q(n_2639));
   AOI211_X2_50_SVT g78581__7482 (.A0(DPATH_RF_MEMORY_18__4_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2441),
	.C0(n_2569),
	.Q(n_2638));
   AOI211_X2_50_SVT g78582__4733 (.A0(DPATH_RF_MEMORY_18__2_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2435),
	.C0(n_2567),
	.Q(n_2637));
   AOI211_X2_50_SVT g78583__6161 (.A0(DPATH_RF_MEMORY_18__1_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2431),
	.C0(n_2566),
	.Q(n_2636));
   AOI211_X2_50_SVT g78584__9315 (.A0(DPATH_RF_MEMORY_18__25_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2426),
	.C0(n_2563),
	.Q(n_2635));
   AOI211_X1_50_SVT g78585__9945 (.A0(DPATH_RF_MEMORY_18__5_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2429),
	.C0(n_2565),
	.Q(n_2634));
   AOI211_X1_50_SVT g78586__2883 (.A0(DPATH_RF_MEMORY_17__18_),
	.A1(n_1414),
	.B0(n_2424),
	.C0(n_2564),
	.Q(n_2633));
   AOI211_X1_50_SVT g78587__2346 (.A0(DPATH_RF_MEMORY_17__17_),
	.A1(n_1414),
	.B0(n_2415),
	.C0(n_2562),
	.Q(n_2632));
   AOI211_X2_50_SVT g78588__1666 (.A0(DPATH_RF_MEMORY_18__25_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2377),
	.C0(n_2561),
	.Q(n_2631));
   AOI211_X2_50_SVT g78589__7410 (.A0(DPATH_RF_MEMORY_18__24_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2374),
	.C0(n_2560),
	.Q(n_2630));
   AOI211_X2_50_SVT g78590__6417 (.A0(DPATH_RF_MEMORY_18__18_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2353),
	.C0(n_2559),
	.Q(n_2629));
   AOI221_X1_50_SVT g78591__5477 (.A0(DPATH_RF_MEMORY_20__21_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__21_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2557),
	.Q(n_2628));
   AOI221_X1_50_SVT g78592__2398 (.A0(DPATH_RF_MEMORY_20__14_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__14_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2558),
	.Q(n_2627));
   AOI221_X1_50_SVT g78593__5107 (.A0(DPATH_RF_MEMORY_20__8_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_19__8_),
	.B1(n_1440),
	.C0(n_2556),
	.Q(n_2626));
   AOI221_X1_50_SVT g78594__6260 (.A0(DPATH_RF_MEMORY_20__7_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_19__7_),
	.B1(n_1440),
	.C0(n_2555),
	.Q(n_2625));
   AOI221_X1_50_SVT g78595__4319 (.A0(DPATH_RF_MEMORY_18__29_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__29_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2573),
	.Q(n_2624));
   AOI221_X1_50_SVT g78596__8428 (.A0(DPATH_RF_MEMORY_17__6_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__6_),
	.B1(n_1386),
	.C0(n_2554),
	.Q(n_2623));
   AOI221_X1_50_SVT g78597__5526 (.A0(DPATH_RF_MEMORY_20__7_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__7_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2553),
	.Q(n_2622));
   AOI221_X1_50_SVT g78598__6783 (.A0(DPATH_RF_MEMORY_17__3_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__3_),
	.B1(n_1386),
	.C0(n_2551),
	.Q(n_2621));
   AOI221_X1_50_SVT g78599__3680 (.A0(DPATH_RF_MEMORY_20__6_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__6_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2550),
	.Q(n_2620));
   AOI221_X0_50_SVT g78600__1617 (.A0(DPATH_RF_MEMORY_21__0_),
	.A1(n_1436),
	.B0(DPATH_RF_MEMORY_22__0_),
	.B1(FE_OFN65_n_1438),
	.C0(n_2549),
	.Q(n_2619));
   AOI221_X1_50_SVT g78601__2802 (.A0(DPATH_RF_MEMORY_20__3_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__3_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2548),
	.Q(n_2618));
   AOI221_X1_50_SVT g78602__1705 (.A0(DPATH_RF_MEMORY_20__2_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__2_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2547),
	.Q(n_2617));
   AOI221_X1_50_SVT g78603__5122 (.A0(DPATH_RF_MEMORY_17__24_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__24_),
	.B1(FE_OFN35_n_1385),
	.C0(n_2546),
	.Q(n_2616));
   AOI221_X1_50_SVT g78604__8246 (.A0(DPATH_RF_MEMORY_17__30_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__30_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2545),
	.Q(n_2615));
   AOI221_X1_50_SVT g78605__7098 (.A0(DPATH_RF_MEMORY_17__29_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__29_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2544),
	.Q(n_2614));
   AOI221_X1_50_SVT g78606__6131 (.A0(DPATH_RF_MEMORY_17__26_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__26_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2543),
	.Q(n_2613));
   AOI221_X1_50_SVT g78607__1881 (.A0(DPATH_RF_MEMORY_20__30_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__30_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2542),
	.Q(n_2612));
   AOI221_X1_50_SVT g78608__5115 (.A0(DPATH_RF_MEMORY_20__13_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__13_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2541),
	.Q(n_2611));
   AOI221_X1_50_SVT g78609__7482 (.A0(DPATH_RF_MEMORY_17__23_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__23_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2540),
	.Q(n_2610));
   AOI221_X1_50_SVT g78610__4733 (.A0(DPATH_RF_MEMORY_21__22_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__22_),
	.B1(FE_OFN65_n_1438),
	.C0(n_2539),
	.Q(n_2609));
   AOI221_X1_50_SVT g78611__6161 (.A0(DPATH_RF_MEMORY_20__21_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__21_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2538),
	.Q(n_2608));
   AOI221_X1_50_SVT g78612__9315 (.A0(DPATH_RF_MEMORY_20__22_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__22_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2537),
	.Q(n_2607));
   AOI221_X1_50_SVT g78613__9945 (.A0(DPATH_RF_MEMORY_20__17_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__17_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2536),
	.Q(n_2606));
   AOI221_X1_50_SVT g78614__2883 (.A0(DPATH_RF_MEMORY_20__16_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__16_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2535),
	.Q(n_2605));
   AOI221_X1_50_SVT g78615__2346 (.A0(DPATH_RF_MEMORY_17__15_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__15_),
	.B1(FE_OFN36_n_1386),
	.C0(n_2534),
	.Q(n_2604));
   AOI211_X2_50_SVT g78616__1666 (.A0(DPATH_RF_MEMORY_20__12_),
	.A1(FE_OFN52_n_1408),
	.B0(n_2164),
	.C0(n_2471),
	.Q(n_2603));
   AOI221_X1_50_SVT g78617__7410 (.A0(DPATH_RF_MEMORY_20__20_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_21__20_),
	.B1(n_1424),
	.C0(n_2531),
	.Q(n_2602));
   INV_A_OAI211_X2_50_SVT g78618__6417 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__19_),
	.B0(n_2356),
	.C0(n_2355),
	.Q(n_2601));
   AOI221_X1_50_SVT g78619__5477 (.A0(DPATH_RF_MEMORY_20__23_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_21__23_),
	.B1(n_1424),
	.C0(n_2509),
	.Q(n_2600));
   AOI221_X1_50_SVT g78620__2398 (.A0(DPATH_RF_MEMORY_20__28_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_21__28_),
	.B1(FE_OFN64_n_1436),
	.C0(n_2506),
	.Q(n_2599));
   AOI221_X1_50_SVT g78621__5107 (.A0(DPATH_RF_MEMORY_22__27_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_19__27_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2504),
	.Q(n_2598));
   AOI221_X1_50_SVT g78622__6260 (.A0(DPATH_RF_MEMORY_20__20_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_21__20_),
	.B1(FE_OFN64_n_1436),
	.C0(n_2496),
	.Q(n_2597));
   AOI221_X1_50_SVT g78623__4319 (.A0(DPATH_RF_MEMORY_22__19_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_19__19_),
	.B1(FE_OFN66_n_1440),
	.C0(n_2493),
	.Q(n_2596));
   AOI221_X1_50_SVT g78624__8428 (.A0(DPATH_RF_MEMORY_19__31_),
	.A1(FE_OFN44_n_1396),
	.B0(DPATH_RF_MEMORY_22__31_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2518),
	.Q(n_2595));
   AOI221_X0_50_SVT g78625__5526 (.A0(DPATH_RF_MEMORY_21__4_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_19__4_),
	.B1(FE_OFN44_n_1396),
	.C0(n_2520),
	.Q(n_2594));
   AOI221_X0_50_SVT g78626__6783 (.A0(DPATH_RF_MEMORY_21__9_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__9_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2532),
	.Q(n_2593));
   INV_A_OAI211_X1_50_SVT g78627__3680 (.A0(n_1384),
	.A1N(DPATH_RF_MEMORY_31__26_),
	.B0(n_2465),
	.C0(n_2151),
	.Q(n_2592));
   AOI221_X0_50_SVT g78628__1617 (.A0(DPATH_RF_MEMORY_21__8_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__8_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2529),
	.Q(n_2591));
   AOI221_X0_50_SVT g78629__2802 (.A0(DPATH_RF_MEMORY_21__28_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__28_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2516),
	.Q(n_2590));
   AOI221_X1_50_SVT g78630__1705 (.A0(DPATH_RF_MEMORY_21__1_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__1_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2514),
	.Q(n_2589));
   AOI221_X0_50_SVT g78631__5122 (.A0(DPATH_RF_MEMORY_21__16_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__16_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2513),
	.Q(n_2588));
   AOI221_X1_50_SVT g78632__8246 (.A0(DPATH_RF_MEMORY_21__31_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__31_),
	.B1(FE_OFN65_n_1438),
	.C0(n_2511),
	.Q(n_2587));
   AOI221_X0_50_SVT g78633__7098 (.A0(DPATH_RF_MEMORY_21__14_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__14_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2505),
	.Q(n_2586));
   AOI221_X0_50_SVT g78634__6131 (.A0(DPATH_RF_MEMORY_21__27_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__27_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2500),
	.Q(n_2585));
   AOI221_X0_50_SVT g78635__1881 (.A0(DPATH_RF_MEMORY_21__11_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__11_),
	.B1(FE_OFN25_n_1331),
	.C0(n_2492),
	.Q(n_2584));
   INV_A_OAI211_X1_50_SVT g78636__5115 (.A0(FE_OFN56_n_1415),
	.A1N(DPATH_RF_MEMORY_17__31_),
	.B0(n_2417),
	.C0(n_2360),
	.Q(n_2583));
   INV_A_OAI211_X2_50_SVT g78637__7482 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__12_),
	.B0(n_2470),
	.C0(n_2469),
	.Q(n_2582));
   INV_A_OAI211_X2_50_SVT g78638__4733 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__10_),
	.B0(n_2460),
	.C0(n_2461),
	.Q(n_2581));
   INV_A_OAI211_X1_50_SVT g78639__6161 (.A0(n_1418),
	.A1N(DPATH_RF_MEMORY_18__20_),
	.B0(n_2456),
	.C0(n_2452),
	.Q(n_2580));
   INV_A_OAI211_X1_50_SVT g78640__9315 (.A0(n_1419),
	.A1N(DPATH_RF_MEMORY_18__4_),
	.B0(n_2421),
	.C0(n_2422),
	.Q(n_2579));
   INV_A_OAI211_X2_50_SVT g78641__9945 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__28_),
	.B0(n_2389),
	.C0(n_2388),
	.Q(n_2578));
   INV_A_OAI211_X1_50_SVT g78642__2883 (.A0(n_1419),
	.A1N(DPATH_RF_MEMORY_18__23_),
	.B0(n_2384),
	.C0(n_2378),
	.Q(n_2577));
   INV_A_OAI211_X2_50_SVT g78643__2346 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__27_),
	.B0(n_2383),
	.C0(n_2385),
	.Q(n_2576));
   INV_A_OAI211_X2_50_SVT g78644__1666 (.A0(n_1431),
	.A1N(DPATH_RF_MEMORY_18__20_),
	.B0(n_2359),
	.C0(n_2358),
	.Q(n_2575));
   AOI221_X1_50_SVT g78645__7410 (.A0(DPATH_RF_MEMORY_20__10_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_21__10_),
	.B1(n_1436),
	.C0(n_2487),
	.Q(n_2574));
   NAND4_X1_50_SVT g78646__6417 (.A(n_2123),
	.B(n_1980),
	.C(n_1934),
	.D(n_2244),
	.Q(n_2573));
   NAND4_X2_50_SVT g78647__5477 (.A(n_2463),
	.B(n_2259),
	.C(n_1494),
	.D(n_2139),
	.Q(n_2572));
   NAND4_X2_50_SVT g78648__2398 (.A(n_2457),
	.B(n_2258),
	.C(n_2013),
	.D(n_2097),
	.Q(n_2571));
   NAND4_X2_50_SVT g78649__5107 (.A(n_2443),
	.B(n_2253),
	.C(n_2021),
	.D(n_2020),
	.Q(n_2570));
   NAND4_X2_50_SVT g78650__6260 (.A(n_2439),
	.B(n_2252),
	.C(n_2002),
	.D(n_2001),
	.Q(n_2569));
   NAND4T_X0_50_SVT g78651__4319 (.A(n_2432),
	.B(n_2250),
	.C(n_1973),
	.D(n_1979),
	.Q(n_2568));
   NAND4_X2_50_SVT g78652__8428 (.A(n_2433),
	.B(n_2249),
	.C(n_1972),
	.D(n_1971),
	.Q(n_2567));
   NAND4_X2_50_SVT g78653__5526 (.A(n_2430),
	.B(n_2247),
	.C(n_1958),
	.D(n_1957),
	.Q(n_2566));
   NAND4T_X0_50_SVT g78654__6783 (.A(n_2425),
	.B(n_2245),
	.C(n_1933),
	.D(n_1938),
	.Q(n_2565));
   NAND4T_X0_50_SVT g78655__3680 (.A(n_2420),
	.B(n_2243),
	.C(n_1907),
	.D(n_1912),
	.Q(n_2564));
   NAND4_X1_50_SVT g78656__1617 (.A(n_1906),
	.B(n_2242),
	.C(n_1900),
	.D(n_2416),
	.Q(n_2563));
   NAND4T_X0_50_SVT g78657__2802 (.A(n_2409),
	.B(n_2240),
	.C(n_1862),
	.D(n_1860),
	.Q(n_2562));
   NAND4_X2_50_SVT g78658__1705 (.A(n_2376),
	.B(n_2232),
	.C(n_1670),
	.D(n_1669),
	.Q(n_2561));
   NAND4_X2_50_SVT g78659__5122 (.A(n_2373),
	.B(n_2231),
	.C(n_1655),
	.D(n_1656),
	.Q(n_2560));
   NAND4_X2_50_SVT g78660__8246 (.A(n_2351),
	.B(n_2223),
	.C(n_1540),
	.D(n_1539),
	.Q(n_2559));
   NAND4T_X0_50_SVT g78661__7098 (.A(n_2233),
	.B(n_2187),
	.C(n_2189),
	.D(n_2186),
	.Q(n_2558));
   NAND4_X2_50_SVT g78662__6131 (.A(n_2260),
	.B(n_2183),
	.C(n_2177),
	.D(n_2168),
	.Q(n_2557));
   NAND4T_X0_50_SVT g78663__1881 (.A(n_2257),
	.B(n_2078),
	.C(n_2079),
	.D(n_2076),
	.Q(n_2556));
   NAND4T_X0_50_SVT g78664__5115 (.A(n_2256),
	.B(n_2058),
	.C(n_2060),
	.D(n_2056),
	.Q(n_2555));
   NAND4T_X0_50_SVT g78665__7482 (.A(n_2255),
	.B(n_2035),
	.C(n_2037),
	.D(n_2038),
	.Q(n_2554));
   NAND4_X1_50_SVT g78666__4733 (.A(n_2025),
	.B(n_2031),
	.C(n_2026),
	.D(n_2254),
	.Q(n_2553));
   NAND4_X2_50_SVT g78667__6161 (.A(n_2473),
	.B(n_2261),
	.C(n_2169),
	.D(n_2167),
	.Q(n_2552));
   NAND4T_X0_50_SVT g78668__9315 (.A(n_2251),
	.B(n_2016),
	.C(n_1985),
	.D(n_1984),
	.Q(n_2551));
   NAND4_X2_50_SVT g78669__9945 (.A(n_2248),
	.B(n_1977),
	.C(n_1475),
	.D(n_1870),
	.Q(n_2550));
   NAND4T_X0_50_SVT g78670__2883 (.A(n_2246),
	.B(n_1936),
	.C(n_1935),
	.D(n_1937),
	.Q(n_2549));
   NAND4_X2_50_SVT g78671__2346 (.A(n_2241),
	.B(n_1882),
	.C(n_1883),
	.D(n_1884),
	.Q(n_2548));
   NAND4_X1_50_SVT g78672__1666 (.A(n_1858),
	.B(n_1861),
	.C(n_1859),
	.D(n_2239),
	.Q(n_2547));
   NAND4_X1_50_SVT g78673__7410 (.A(n_1785),
	.B(n_1796),
	.C(n_1792),
	.D(n_2236),
	.Q(n_2546));
   NAND4T_X0_50_SVT g78674__6417 (.A(n_2235),
	.B(n_1766),
	.C(n_1767),
	.D(n_1763),
	.Q(n_2545));
   NAND4T_X0_50_SVT g78675__5477 (.A(n_2234),
	.B(n_1747),
	.C(n_1748),
	.D(n_1745),
	.Q(n_2544));
   NAND4T_X0_50_SVT g78676__2398 (.A(n_2262),
	.B(n_1688),
	.C(n_1687),
	.D(n_1689),
	.Q(n_2543));
   NAND4T_X0_50_SVT g78677__5107 (.A(n_2225),
	.B(n_1679),
	.C(n_1651),
	.D(n_1700),
	.Q(n_2542));
   NAND4_X1_50_SVT g78678__6260 (.A(n_1643),
	.B(n_1647),
	.C(n_1638),
	.D(n_2230),
	.Q(n_2541));
   NAND4T_X0_50_SVT g78679__4319 (.A(n_2229),
	.B(n_1632),
	.C(n_1635),
	.D(n_1634),
	.Q(n_2540));
   NAND4T_X0_50_SVT g78680__8428 (.A(n_2227),
	.B(n_1612),
	.C(n_1613),
	.D(n_1611),
	.Q(n_2539));
   NAND4T_X0_50_SVT g78681__5526 (.A(n_2226),
	.B(n_1591),
	.C(n_1593),
	.D(n_1594),
	.Q(n_2538));
   NAND4_X1_50_SVT g78682__6783 (.A(n_1560),
	.B(n_1571),
	.C(n_1566),
	.D(n_2224),
	.Q(n_2537));
   NAND4T_X0_50_SVT g78683__3680 (.A(n_2222),
	.B(n_1519),
	.C(n_1522),
	.D(n_1520),
	.Q(n_2536));
   NAND4T_X0_50_SVT g78684__1617 (.A(n_2220),
	.B(n_1498),
	.C(n_1501),
	.D(n_1499),
	.Q(n_2535));
   NAND4T_X0_50_SVT g78685__2802 (.A(n_2219),
	.B(n_1474),
	.C(n_1478),
	.D(n_1476),
	.Q(n_2534));
   AOI21_X1_50_SVT g78686__1705 (.A0(DPATH_RF_MEMORY_17__10_),
	.A1(n_1415),
	.B0(n_2476),
	.Q(n_2533));
   AO21_X2_50_SVT g78687__5122 (.A0(DPATH_RF_MEMORY_31__9_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2472),
	.Q(n_2532));
   AO21_X2_50_SVT g78688__8246 (.A0(DPATH_RF_MEMORY_19__20_),
	.A1(FE_OFN44_n_1396),
	.B0(n_2464),
	.Q(n_2531));
   AOI21_X2_50_SVT g78689__7098 (.A0(DPATH_RF_MEMORY_18__14_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2339),
	.Q(n_2530));
   AO21_X2_50_SVT g78690__6131 (.A0(DPATH_RF_MEMORY_31__8_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2459),
	.Q(n_2529));
   AOI21_X2_50_SVT g78691__1881 (.A0(DPATH_RF_MEMORY_18__8_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2454),
	.Q(n_2528));
   AOI21_X2_50_SVT g78692__5115 (.A0(DPATH_RF_MEMORY_17__7_),
	.A1(n_1415),
	.B0(n_2450),
	.Q(n_2527));
   AOI21_X2_50_SVT g78693__7482 (.A0(DPATH_RF_MEMORY_18__7_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2451),
	.Q(n_2526));
   AOI21_X2_50_SVT g78694__4733 (.A0(DPATH_RF_MEMORY_18__6_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2447),
	.Q(n_2525));
   AOI21_X1_50_SVT g78695__6161 (.A0(DPATH_RF_MEMORY_17__30_),
	.A1(n_1414),
	.B0(n_2434),
	.Q(n_2524));
   AOI21_X0_50_SVT g78696__9315 (.A0(DPATH_RF_MEMORY_18__6_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2440),
	.Q(n_2523));
   AOI21_X2_50_SVT g78697__9945 (.A0(DPATH_RF_MEMORY_18__3_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2437),
	.Q(n_2522));
   AOI21_X2_50_SVT g78698__2883 (.A0(DPATH_RF_MEMORY_18__0_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2428),
	.Q(n_2521));
   AO21_X2_50_SVT g78699__2346 (.A0(DPATH_RF_MEMORY_20__4_),
	.A1(FE_OFN41_n_1392),
	.B0(n_2423),
	.Q(n_2520));
   AOI21_X1_50_SVT g78700__1666 (.A0(DPATH_RF_MEMORY_18__3_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2419),
	.Q(n_2519));
   AO21_X2_50_SVT g78701__7410 (.A0(DPATH_RF_MEMORY_20__31_),
	.A1(FE_OFN41_n_1392),
	.B0(n_2394),
	.Q(n_2518));
   AOI21_X1_50_SVT g78702__6417 (.A0(DPATH_RF_MEMORY_17__2_),
	.A1(n_1415),
	.B0(n_2414),
	.Q(n_2517));
   AO21_X2_50_SVT g78703__5477 (.A0(DPATH_RF_MEMORY_31__28_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2402),
	.Q(n_2516));
   AOI21_X2_50_SVT g78704__2398 (.A0(DPATH_RF_MEMORY_18__24_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2411),
	.Q(n_2515));
   AO21_X2_50_SVT g78705__5107 (.A0(DPATH_RF_MEMORY_31__1_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2410),
	.Q(n_2514));
   AO21_X2_50_SVT g78706__6260 (.A0(DPATH_RF_MEMORY_31__16_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2406),
	.Q(n_2513));
   AOI21_X2_50_SVT g78707__4319 (.A0(DPATH_RF_MEMORY_17__0_),
	.A1(n_1415),
	.B0(n_2404),
	.Q(n_2512));
   AO21_X2_50_SVT g78708__8428 (.A0(DPATH_RF_MEMORY_31__31_),
	.A1(FE_OFN36_n_1386),
	.B0(n_2401),
	.Q(n_2511));
   AOI21_X2_50_SVT g78709__5526 (.A0(DPATH_RF_MEMORY_18__30_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2399),
	.Q(n_2510));
   AO21_X2_50_SVT g78710__6783 (.A0(DPATH_RF_MEMORY_19__23_),
	.A1(FE_OFN44_n_1396),
	.B0(n_2393),
	.Q(n_2509));
   AOI21_X1_50_SVT g78711__3680 (.A0(DPATH_RF_MEMORY_17__15_),
	.A1(n_1414),
	.B0(n_2392),
	.Q(n_2508));
   AOI21_X2_50_SVT g78712__1617 (.A0(DPATH_RF_MEMORY_18__29_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2395),
	.Q(n_2507));
   AO21_X2_50_SVT g78713__2802 (.A0(DPATH_RF_MEMORY_19__28_),
	.A1(FE_OFN66_n_1440),
	.B0(n_2390),
	.Q(n_2506));
   AO21_X2_50_SVT g78714__1705 (.A0(DPATH_RF_MEMORY_31__14_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2387),
	.Q(n_2505));
   AO21_X2_50_SVT g78715__5122 (.A0(DPATH_RF_MEMORY_21__27_),
	.A1(FE_OFN64_n_1436),
	.B0(n_2386),
	.Q(n_2504));
   AOI21_X2_50_SVT g78716__8246 (.A0(DPATH_RF_MEMORY_18__26_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2382),
	.Q(n_2503));
   AOI21_X2_50_SVT g78717__7098 (.A0(DPATH_RF_MEMORY_17__13_),
	.A1(n_1415),
	.B0(n_2379),
	.Q(n_2502));
   AOI21_X1_50_SVT g78718__6131 (.A0(DPATH_RF_MEMORY_18__22_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2371),
	.Q(n_2501));
   AO21_X2_50_SVT g78719__1881 (.A0(DPATH_RF_MEMORY_31__27_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2370),
	.Q(n_2500));
   AOI21_X2_50_SVT g78720__5115 (.A0(DPATH_RF_MEMORY_18__23_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2372),
	.Q(n_2499));
   AOI21_X2_50_SVT g78721__7482 (.A0(DPATH_RF_MEMORY_18__22_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2367),
	.Q(n_2498));
   AOI21_X2_50_SVT g78722__4733 (.A0(DPATH_RF_MEMORY_18__21_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2365),
	.Q(n_2497));
   AO21_X2_50_SVT g78723__6161 (.A0(DPATH_RF_MEMORY_19__20_),
	.A1(FE_OFN66_n_1440),
	.B0(n_2362),
	.Q(n_2496));
   AOI21_X1_50_SVT g78724__9315 (.A0(DPATH_RF_MEMORY_17__12_),
	.A1(n_1414),
	.B0(n_2361),
	.Q(n_2495));
   AOI21_X2_50_SVT g78725__9945 (.A0(DPATH_RF_MEMORY_17__29_),
	.A1(n_1414),
	.B0(n_2352),
	.Q(n_2494));
   AO21_X2_50_SVT g78726__2883 (.A0(DPATH_RF_MEMORY_21__19_),
	.A1(FE_OFN64_n_1436),
	.B0(n_2357),
	.Q(n_2493));
   AO21_X2_50_SVT g78727__2346 (.A0(DPATH_RF_MEMORY_31__11_),
	.A1(FE_OFN35_n_1385),
	.B0(n_2354),
	.Q(n_2492));
   AOI21_X2_50_SVT g78728__1666 (.A0(DPATH_RF_MEMORY_18__21_),
	.A1(FE_OFN57_n_1419),
	.B0(n_2349),
	.Q(n_2491));
   AOI21_X2_50_SVT g78729__7410 (.A0(DPATH_RF_MEMORY_18__17_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2347),
	.Q(n_2490));
   AOI21_X2_50_SVT g78730__6417 (.A0(DPATH_RF_MEMORY_18__16_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2345),
	.Q(n_2489));
   AOI21_X2_50_SVT g78731__5477 (.A0(DPATH_RF_MEMORY_18__15_),
	.A1(FE_OFN63_n_1432),
	.B0(n_2342),
	.Q(n_2488));
   AO21_X2_50_SVT g78732__2398 (.A0(DPATH_RF_MEMORY_22__10_),
	.A1(n_1438),
	.B0(n_2462),
	.Q(n_2487));
   AOI221_X1_50_SVT g78733__5107 (.A0(DPATH_RF_MEMORY_1__7_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__7_),
	.B1(n_1434),
	.C0(n_2326),
	.Q(n_2486));
   AOI221_X0_50_SVT g78734__6260 (.A0(DPATH_RF_MEMORY_13__8_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__8_),
	.B1(n_1412),
	.C0(n_2271),
	.Q(n_2485));
   AOI221_X0_50_SVT g78735__4319 (.A0(DPATH_RF_MEMORY_13__26_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__26_),
	.B1(n_1412),
	.C0(n_2270),
	.Q(n_2484));
   AOI221_X1_50_SVT g78736__8428 (.A0(DPATH_RF_MEMORY_8__1_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__1_),
	.B1(n_1403),
	.C0(n_2269),
	.Q(n_2483));
   AOI221_X1_50_SVT g78737__5526 (.A0(DPATH_RF_MEMORY_5__16_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__16_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2268),
	.Q(n_2482));
   AOI221_X0_50_SVT g78738__6783 (.A0(DPATH_RF_MEMORY_4__28_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__28_),
	.B1(n_1420),
	.C0(n_2266),
	.Q(n_2481));
   AOI221_X1_50_SVT g78739__3680 (.A0(DPATH_RF_MEMORY_8__31_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__31_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2267),
	.Q(n_2480));
   AOI221_X2_50_SVT g78740__1617 (.A0(DPATH_RF_MEMORY_5__14_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__14_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2265),
	.Q(n_2479));
   AOI221_X1_50_SVT g78741__2802 (.A0(DPATH_RF_MEMORY_12__27_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__27_),
	.B1(FE_OFN40_n_1391),
	.C0(n_2264),
	.Q(n_2478));
   AOI221_X1_50_SVT g78742__1705 (.A0(DPATH_RF_MEMORY_4__11_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__11_),
	.B1(n_1420),
	.C0(n_2263),
	.Q(n_2477));
   NAND4_X2_50_SVT g78743__5122 (.A(n_2197),
	.B(n_2192),
	.C(n_2190),
	.D(n_2184),
	.Q(n_2476));
   AOI221_X1_50_SVT g78744__8246 (.A0(DPATH_RF_MEMORY_29__14_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__14_),
	.B1(n_1378),
	.C0(n_2318),
	.Q(n_2475));
   NAND4T_X0_50_SVT g78745__7098 (.A(n_2178),
	.B(n_2176),
	.C(n_2179),
	.D(n_2175),
	.Q(n_2474));
   AOI221_X1_50_SVT g78746__6131 (.A0(DPATH_RF_MEMORY_24__13_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__13_),
	.B1(n_1445),
	.C0(n_2337),
	.Q(n_2473));
   NAND4_X2_50_SVT g78747__1881 (.A(n_2166),
	.B(n_2159),
	.C(n_2161),
	.D(n_2155),
	.Q(n_2472));
   NAND4T_X0_50_SVT g78748__5115 (.A(n_2157),
	.B(n_2162),
	.C(n_2160),
	.D(n_2158),
	.Q(n_2471));
   AOI221_X1_50_SVT g78749__7482 (.A0(DPATH_RF_MEMORY_9__12_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__12_),
	.B1(n_1399),
	.C0(n_2336),
	.Q(n_2470));
   AOI221_X1_50_SVT g78750__4733 (.A0(DPATH_RF_MEMORY_4__12_),
	.A1(n_1380),
	.B0(DPATH_RF_MEMORY_3__12_),
	.B1(n_1446),
	.C0(n_2335),
	.Q(n_2469));
   AOI221_X1_50_SVT g78751__6161 (.A0(DPATH_RF_MEMORY_8__29_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__29_),
	.B1(n_1403),
	.C0(n_2334),
	.Q(n_2468));
   NAND4T_X0_50_SVT g78752__9315 (.A(n_2140),
	.B(n_2144),
	.C(n_2143),
	.D(n_2141),
	.Q(n_2467));
   NAND4_X2_50_SVT g78753__9945 (.A(n_2137),
	.B(n_2142),
	.C(n_2131),
	.D(n_2135),
	.Q(n_2466));
   AOI221_X0_50_SVT g78754__2883 (.A0(DPATH_RF_MEMORY_28__26_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__26_),
	.B1(FE_OFN55_n_1413),
	.C0(n_2327),
	.Q(n_2465));
   NAND4_X2_50_SVT g78755__2346 (.A(n_2138),
	.B(n_2122),
	.C(n_2133),
	.D(n_2117),
	.Q(n_2464));
   AOI221_X1_50_SVT g78756__1666 (.A0(DPATH_RF_MEMORY_1__11_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__11_),
	.B1(n_1434),
	.C0(n_2333),
	.Q(n_2463));
   NAND4T_X0_50_SVT g78757__7410 (.A(n_2126),
	.B(n_2128),
	.C(n_2125),
	.D(n_2124),
	.Q(n_2462));
   AOI221_X1_50_SVT g78758__6417 (.A0(DPATH_RF_MEMORY_29__10_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__10_),
	.B1(n_1378),
	.C0(n_2332),
	.Q(n_2461));
   AOI221_X1_50_SVT g78759__5477 (.A0(DPATH_RF_MEMORY_8__10_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__10_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2331),
	.Q(n_2460));
   NAND4_X2_50_SVT g78760__2398 (.A(n_2108),
	.B(n_2112),
	.C(n_2105),
	.D(n_2104),
	.Q(n_2459));
   NAND4T_X0_50_SVT g78761__5107 (.A(n_1966),
	.B(n_2103),
	.C(n_2107),
	.D(n_2106),
	.Q(n_2458));
   AOI221_X1_50_SVT g78762__6260 (.A0(DPATH_RF_MEMORY_13__9_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__9_),
	.B1(FE_OFN48_n_1401),
	.C0(n_2330),
	.Q(n_2457));
   AOI221_X0_50_SVT g78763__4319 (.A0(DPATH_RF_MEMORY_25__20_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__20_),
	.B1(FE_OFN53_n_1409),
	.C0(n_2329),
	.Q(n_2456));
   NAND4_X2_50_SVT g78764__8428 (.A(n_2085),
	.B(n_1510),
	.C(n_2080),
	.D(n_2072),
	.Q(n_2455));
   NAND4_X2_50_SVT g78765__5526 (.A(n_2093),
	.B(n_2092),
	.C(n_2090),
	.D(n_2089),
	.Q(n_2454));
   AOI221_X1_50_SVT g78766__6783 (.A0(DPATH_RF_MEMORY_25__8_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__8_),
	.B1(FE_OFN38_n_1389),
	.C0(n_2328),
	.Q(n_2453));
   AOI221_X1_50_SVT g78767__3680 (.A0(DPATH_RF_MEMORY_1__20_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__20_),
	.B1(n_1427),
	.C0(n_2325),
	.Q(n_2452));
   NAND4T_X0_50_SVT g78768__1617 (.A(n_2073),
	.B(n_2071),
	.C(n_2074),
	.D(n_2070),
	.Q(n_2451));
   NAND4_X2_50_SVT g78769__2802 (.A(n_2062),
	.B(n_2068),
	.C(n_2061),
	.D(n_2057),
	.Q(n_2450));
   AOI221_X0_50_SVT g78770__1705 (.A0(DPATH_RF_MEMORY_12__9_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__9_),
	.B1(FE_OFN40_n_1391),
	.C0(n_2272),
	.Q(n_2449));
   AOI221_X0_50_SVT g78771__5122 (.A0(DPATH_RF_MEMORY_24__7_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__7_),
	.B1(FE_OFN33_n_1381),
	.C0(n_2324),
	.Q(n_2448));
   NAND4T_X0_50_SVT g78772__8246 (.A(n_2050),
	.B(n_2048),
	.C(n_2052),
	.D(n_2051),
	.Q(n_2447));
   AOI221_X1_50_SVT g78773__7098 (.A0(DPATH_RF_MEMORY_4__6_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__6_),
	.B1(n_1446),
	.C0(n_2323),
	.Q(n_2446));
   AOI221_X1_50_SVT g78774__6131 (.A0(DPATH_RF_MEMORY_4__26_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__26_),
	.B1(n_1420),
	.C0(n_2321),
	.Q(n_2445));
   NAND4T_X0_50_SVT g78775__1881 (.A(n_2028),
	.B(n_2027),
	.C(n_2029),
	.D(n_2030),
	.Q(n_2444));
   AOI221_X1_50_SVT g78776__5115 (.A0(DPATH_RF_MEMORY_29__5_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__5_),
	.B1(n_1378),
	.C0(n_2322),
	.Q(n_2443));
   NAND4_X2_50_SVT g78777__7482 (.A(n_2015),
	.B(n_1999),
	.C(n_2009),
	.D(n_1991),
	.Q(n_2442));
   NAND4T_X0_50_SVT g78778__4733 (.A(n_1921),
	.B(n_2014),
	.C(n_2010),
	.D(n_1910),
	.Q(n_2441));
   NAND4_X2_50_SVT g78779__6161 (.A(n_2011),
	.B(n_2008),
	.C(n_2003),
	.D(n_2006),
	.Q(n_2440));
   AOI221_X1_50_SVT g78780__9315 (.A0(DPATH_RF_MEMORY_29__4_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__4_),
	.B1(n_1378),
	.C0(n_2320),
	.Q(n_2439));
   AOI221_X1_50_SVT g78781__9945 (.A0(DPATH_RF_MEMORY_4__6_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__6_),
	.B1(n_1420),
	.C0(n_2319),
	.Q(n_2438));
   NAND4_X2_50_SVT g78782__2883 (.A(n_1997),
	.B(n_1996),
	.C(n_1995),
	.D(n_1994),
	.Q(n_2437));
   AOI221_X1_50_SVT g78783__2346 (.A0(DPATH_RF_MEMORY_29__3_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__3_),
	.B1(n_1378),
	.C0(n_2338),
	.Q(n_2436));
   NAND4T_X0_50_SVT g78784__1666 (.A(n_1975),
	.B(n_1976),
	.C(n_1551),
	.D(n_1974),
	.Q(n_2435));
   NAND4_X2_50_SVT g78785__7410 (.A(n_1930),
	.B(n_1983),
	.C(n_1909),
	.D(n_1888),
	.Q(n_2434));
   AOI221_X1_50_SVT g78786__6417 (.A0(DPATH_RF_MEMORY_1__2_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__2_),
	.B1(n_1434),
	.C0(n_2317),
	.Q(n_2433));
   AOI221_X1_50_SVT g78787__5477 (.A0(DPATH_RF_MEMORY_4__19_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__19_),
	.B1(n_1420),
	.C0(n_2315),
	.Q(n_2432));
   NAND4T_X0_50_SVT g78788__2398 (.A(n_1960),
	.B(n_1959),
	.C(n_1961),
	.D(n_1592),
	.Q(n_2431));
   AOI221_X1_50_SVT g78789__5107 (.A0(DPATH_RF_MEMORY_1__1_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__1_),
	.B1(n_1434),
	.C0(n_2316),
	.Q(n_2430));
   NAND4_X2_50_SVT g78790__6260 (.A(n_1954),
	.B(n_1946),
	.C(n_1951),
	.D(n_1943),
	.Q(n_2429));
   NAND4_X2_50_SVT g78791__4319 (.A(n_1950),
	.B(n_1949),
	.C(n_1947),
	.D(n_1945),
	.Q(n_2428));
   AOI221_X1_50_SVT g78792__8428 (.A0(DPATH_RF_MEMORY_24__0_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__0_),
	.B1(n_1445),
	.C0(n_2314),
	.Q(n_2427));
   NAND4_X2_50_SVT g78793__5526 (.A(n_1931),
	.B(n_1926),
	.C(n_1914),
	.D(n_1923),
	.Q(n_2426));
   AOI221_X1_50_SVT g78794__6783 (.A0(DPATH_RF_MEMORY_5__5_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__5_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2313),
	.Q(n_2425));
   NAND4_X2_50_SVT g78795__3680 (.A(n_2129),
	.B(n_1919),
	.C(n_1915),
	.D(n_1922),
	.Q(n_2424));
   NAND4_X2_50_SVT g78796__1617 (.A(n_1924),
	.B(n_1917),
	.C(n_1918),
	.D(n_1916),
	.Q(n_2423));
   AOI221_X1_50_SVT g78797__2802 (.A0(DPATH_RF_MEMORY_9__4_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__4_),
	.B1(n_1417),
	.C0(n_2312),
	.Q(n_2422));
   AOI221_X1_50_SVT g78798__1705 (.A0(DPATH_RF_MEMORY_5__4_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__4_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2311),
	.Q(n_2421));
   AOI221_X1_50_SVT g78799__5122 (.A0(DPATH_RF_MEMORY_8__18_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__18_),
	.B1(n_1403),
	.C0(n_2310),
	.Q(n_2420));
   NAND4_X2_50_SVT g78800__8246 (.A(n_1901),
	.B(n_1898),
	.C(n_1899),
	.D(n_1895),
	.Q(n_2419));
   AOI221_X2_50_SVT g78801__7098 (.A0(DPATH_RF_MEMORY_5__3_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__3_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2309),
	.Q(n_2418));
   AOI221_X1_50_SVT g78802__6131 (.A0(DPATH_RF_MEMORY_28__31_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__31_),
	.B1(FE_OFN55_n_1413),
	.C0(n_2304),
	.Q(n_2417));
   AOI221_X1_50_SVT g78803__1881 (.A0(DPATH_RF_MEMORY_4__25_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__25_),
	.B1(n_1420),
	.C0(n_2308),
	.Q(n_2416));
   NAND4_X2_50_SVT g78804__5115 (.A(n_1878),
	.B(n_1871),
	.C(n_1876),
	.D(n_1869),
	.Q(n_2415));
   NAND4_X2_50_SVT g78805__7482 (.A(n_1877),
	.B(n_1875),
	.C(n_1874),
	.D(n_1873),
	.Q(n_2414));
   AOI221_X1_50_SVT g78806__4733 (.A0(DPATH_RF_MEMORY_5__2_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__2_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2307),
	.Q(n_2413));
   AOI221_X1_50_SVT g78807__6161 (.A0(DPATH_RF_MEMORY_24__13_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__13_),
	.B1(FE_OFN33_n_1381),
	.C0(n_2290),
	.Q(n_2412));
   NAND4_X2_50_SVT g78808__9315 (.A(n_1851),
	.B(n_1855),
	.C(n_1846),
	.D(n_1841),
	.Q(n_2411));
   NAND4_X2_50_SVT g78809__9945 (.A(n_1849),
	.B(n_1845),
	.C(n_1847),
	.D(n_1844),
	.Q(n_2410));
   AOI221_X1_50_SVT g78810__2883 (.A0(DPATH_RF_MEMORY_4__17_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__17_),
	.B1(n_1420),
	.C0(n_2305),
	.Q(n_2409));
   AOI221_X1_50_SVT g78811__2346 (.A0(DPATH_RF_MEMORY_25__24_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__24_),
	.B1(FE_OFN53_n_1409),
	.C0(n_2303),
	.Q(n_2408));
   NAND4_X2_50_SVT g78812__1666 (.A(n_1835),
	.B(n_1838),
	.C(n_1834),
	.D(n_1832),
	.Q(n_2407));
   NAND4_X2_50_SVT g78813__7410 (.A(n_1829),
	.B(n_1823),
	.C(n_1825),
	.D(n_1820),
	.Q(n_2406));
   AOI221_X1_50_SVT g78814__6417 (.A0(DPATH_RF_MEMORY_1__0_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__0_),
	.B1(n_1427),
	.C0(n_2302),
	.Q(n_2405));
   NAND4_X2_50_SVT g78815__5477 (.A(n_1814),
	.B(n_1810),
	.C(n_1812),
	.D(n_1808),
	.Q(n_2404));
   NAND4_X2_50_SVT g78816__2398 (.A(n_1803),
	.B(n_1804),
	.C(n_1800),
	.D(n_1798),
	.Q(n_2403));
   NAND4_X2_50_SVT g78817__5107 (.A(n_1837),
	.B(n_1853),
	.C(n_1827),
	.D(n_1813),
	.Q(n_2402));
   NAND4T_X0_50_SVT g78818__6260 (.A(n_1797),
	.B(n_1799),
	.C(n_1794),
	.D(n_1793),
	.Q(n_2401));
   NAND4T_X0_50_SVT g78819__4319 (.A(n_1783),
	.B(n_1784),
	.C(n_1787),
	.D(n_1782),
	.Q(n_2400));
   NAND4T_X0_50_SVT g78820__8428 (.A(n_1777),
	.B(n_1776),
	.C(n_1779),
	.D(n_1778),
	.Q(n_2399));
   AOI221_X1_50_SVT g78821__5526 (.A0(DPATH_RF_MEMORY_5__15_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__15_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2300),
	.Q(n_2398));
   AOI221_X1_50_SVT g78822__6783 (.A0(DPATH_RF_MEMORY_5__30_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__30_),
	.B1(FE_OFN49_n_1404),
	.C0(n_2301),
	.Q(n_2397));
   NAND4_X2_50_SVT g78823__3680 (.A(n_1736),
	.B(n_1755),
	.C(n_1727),
	.D(n_1712),
	.Q(n_2396));
   NAND4_X2_50_SVT g78824__1617 (.A(n_1760),
	.B(n_1759),
	.C(n_1758),
	.D(n_1757),
	.Q(n_2395));
   NAND4T_X0_50_SVT g78825__2802 (.A(n_1886),
	.B(n_1741),
	.C(n_1624),
	.D(n_1615),
	.Q(n_2394));
   NAND4_X2_50_SVT g78826__1705 (.A(n_1746),
	.B(n_1735),
	.C(n_1744),
	.D(n_1731),
	.Q(n_2393));
   NAND4_X2_50_SVT g78827__5122 (.A(n_1751),
	.B(n_1756),
	.C(n_1749),
	.D(n_1743),
	.Q(n_2392));
   AOI221_X1_50_SVT g78828__8246 (.A0(DPATH_RF_MEMORY_29__29_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__29_),
	.B1(n_1378),
	.C0(n_2299),
	.Q(n_2391));
   NAND4T_X0_50_SVT g78829__7098 (.A(n_1733),
	.B(n_1739),
	.C(n_1734),
	.D(n_1737),
	.Q(n_2390));
   AOI221_X1_50_SVT g78830__6131 (.A0(DPATH_RF_MEMORY_13__28_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__28_),
	.B1(FE_OFN48_n_1401),
	.C0(n_2298),
	.Q(n_2389));
   AOI221_X1_50_SVT g78831__1881 (.A0(DPATH_RF_MEMORY_5__28_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__28_),
	.B1(FE_OFN49_n_1404),
	.C0(n_2297),
	.Q(n_2388));
   NAND4_X2_50_SVT g78832__5115 (.A(n_1725),
	.B(n_1719),
	.C(n_1722),
	.D(n_1716),
	.Q(n_2387));
   NAND4T_X0_50_SVT g78833__7482 (.A(n_1720),
	.B(n_1721),
	.C(n_1718),
	.D(n_1717),
	.Q(n_2386));
   AOI221_X1_50_SVT g78834__4733 (.A0(DPATH_RF_MEMORY_28__27_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__27_),
	.B1(FE_OFN31_n_1379),
	.C0(n_2296),
	.Q(n_2385));
   AOI221_X0_50_SVT g78835__6161 (.A0(DPATH_RF_MEMORY_28__23_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__23_),
	.B1(FE_OFN55_n_1413),
	.C0(n_2294),
	.Q(n_2384));
   AOI221_X1_50_SVT g78836__9315 (.A0(DPATH_RF_MEMORY_5__27_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__27_),
	.B1(FE_OFN49_n_1404),
	.C0(n_2295),
	.Q(n_2383));
   NAND4_X2_50_SVT g78837__9945 (.A(n_1706),
	.B(n_1704),
	.C(n_1702),
	.D(n_1703),
	.Q(n_2382));
   NAND4_X2_50_SVT g78838__2883 (.A(n_1699),
	.B(n_1690),
	.C(n_1695),
	.D(n_1686),
	.Q(n_2381));
   AOI221_X1_50_SVT g78839__2346 (.A0(DPATH_RF_MEMORY_29__26_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__26_),
	.B1(n_1378),
	.C0(n_2293),
	.Q(n_2380));
   NAND4_X2_50_SVT g78840__1666 (.A(n_1682),
	.B(n_1677),
	.C(n_1671),
	.D(n_1675),
	.Q(n_2379));
   AOI221_X1_50_SVT g78841__7410 (.A0(DPATH_RF_MEMORY_5__23_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__23_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2291),
	.Q(n_2378));
   NAND4T_X0_50_SVT g78842__6417 (.A(n_1680),
	.B(n_1711),
	.C(n_1681),
	.D(n_1678),
	.Q(n_2377));
   AOI221_X1_50_SVT g78843__5477 (.A0(DPATH_RF_MEMORY_12__25_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__25_),
	.B1(n_1450),
	.C0(n_2292),
	.Q(n_2376));
   AOI221_X1_50_SVT g78844__2398 (.A0(DPATH_RF_MEMORY_4__30_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__30_),
	.B1(n_1420),
	.C0(n_2306),
	.Q(n_2375));
   NAND4T_X0_50_SVT g78845__5107 (.A(n_1661),
	.B(n_1659),
	.C(n_1664),
	.D(n_1663),
	.Q(n_2374));
   AOI221_X1_50_SVT g78846__6260 (.A0(DPATH_RF_MEMORY_1__24_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__24_),
	.B1(n_1434),
	.C0(n_2289),
	.Q(n_2373));
   NAND4T_X0_50_SVT g78847__4319 (.A(n_1645),
	.B(n_1646),
	.C(n_1649),
	.D(n_1644),
	.Q(n_2372));
   NAND4_X2_50_SVT g78848__8428 (.A(n_1648),
	.B(n_1633),
	.C(n_1640),
	.D(n_1628),
	.Q(n_2371));
   NAND4_X2_50_SVT g78849__5526 (.A(n_1637),
	.B(n_1619),
	.C(n_1603),
	.D(n_1579),
	.Q(n_2370));
   AOI221_X1_50_SVT g78850__6783 (.A0(DPATH_RF_MEMORY_8__23_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__23_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2288),
	.Q(n_2369));
   AOI221_X2_50_SVT g78851__3680 (.A0(DPATH_RF_MEMORY_5__22_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__22_),
	.B1(FE_OFN59_n_1423),
	.C0(n_2286),
	.Q(n_2368));
   NAND4_X2_50_SVT g78852__1617 (.A(n_1627),
	.B(n_1625),
	.C(n_1623),
	.D(n_1622),
	.Q(n_2367));
   AOI221_X1_50_SVT g78853__2802 (.A0(DPATH_RF_MEMORY_28__22_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__22_),
	.B1(FE_OFN31_n_1379),
	.C0(n_2287),
	.Q(n_2366));
   NAND4_X2_50_SVT g78854__1705 (.A(n_1608),
	.B(n_1606),
	.C(n_1605),
	.D(n_1604),
	.Q(n_2365));
   AOI221_X1_50_SVT g78855__5122 (.A0(DPATH_RF_MEMORY_4__12_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__12_),
	.B1(n_1420),
	.C0(n_2285),
	.Q(n_2364));
   AOI221_X2_50_SVT g78856__8246 (.A0(DPATH_RF_MEMORY_29__21_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__21_),
	.B1(n_1378),
	.C0(n_2284),
	.Q(n_2363));
   NAND4T_X0_50_SVT g78857__7098 (.A(n_1585),
	.B(n_1584),
	.C(n_1586),
	.D(n_1583),
	.Q(n_2362));
   NAND4_X2_50_SVT g78858__6131 (.A(n_1581),
	.B(n_1582),
	.C(n_1576),
	.D(n_1572),
	.Q(n_2361));
   AOI221_X1_50_SVT g78859__1881 (.A0(DPATH_RF_MEMORY_4__31_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__31_),
	.B1(n_1420),
	.C0(n_2278),
	.Q(n_2360));
   AOI221_X1_50_SVT g78860__5115 (.A0(DPATH_RF_MEMORY_13__20_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__20_),
	.B1(FE_OFN48_n_1401),
	.C0(n_2283),
	.Q(n_2359));
   AOI221_X1_50_SVT g78861__7482 (.A0(DPATH_RF_MEMORY_8__20_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__20_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2282),
	.Q(n_2358));
   NAND4T_X0_50_SVT g78862__4733 (.A(n_1568),
	.B(n_1567),
	.C(n_1569),
	.D(n_1565),
	.Q(n_2357));
   AOI221_X1_50_SVT g78863__6161 (.A0(DPATH_RF_MEMORY_9__19_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__19_),
	.B1(n_1399),
	.C0(n_2281),
	.Q(n_2356));
   AOI221_X1_50_SVT g78864__9315 (.A0(DPATH_RF_MEMORY_1__19_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__19_),
	.B1(n_1434),
	.C0(n_2280),
	.Q(n_2355));
   NAND4_X2_50_SVT g78865__9945 (.A(n_1558),
	.B(n_1552),
	.C(n_1550),
	.D(n_1545),
	.Q(n_2354));
   NAND4T_X0_50_SVT g78866__2883 (.A(n_1548),
	.B(n_1549),
	.C(n_1547),
	.D(n_1546),
	.Q(n_2353));
   NAND4_X2_50_SVT g78867__2346 (.A(n_1538),
	.B(n_1490),
	.C(n_1480),
	.D(n_1836),
	.Q(n_2352));
   AOI221_X1_50_SVT g78868__1666 (.A0(DPATH_RF_MEMORY_29__18_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__18_),
	.B1(n_1378),
	.C0(n_2279),
	.Q(n_2351));
   NAND4_X2_50_SVT g78869__7410 (.A(n_1528),
	.B(n_1509),
	.C(n_1481),
	.D(n_1496),
	.Q(n_2350));
   NAND4_X2_50_SVT g78870__6417 (.A(n_1534),
	.B(n_1518),
	.C(n_1514),
	.D(n_1515),
	.Q(n_2349));
   NAND4_X2_50_SVT g78871__5477 (.A(n_1529),
	.B(n_1524),
	.C(n_1516),
	.D(n_1521),
	.Q(n_2348));
   NAND4_X2_50_SVT g78872__2398 (.A(n_1535),
	.B(n_1533),
	.C(n_1530),
	.D(n_1531),
	.Q(n_2347));
   AOI221_X1_50_SVT g78873__5107 (.A0(DPATH_RF_MEMORY_24__17_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__17_),
	.B1(n_1445),
	.C0(n_2277),
	.Q(n_2346));
   NAND4_X2_50_SVT g78874__6260 (.A(n_1513),
	.B(n_1511),
	.C(n_1507),
	.D(n_1508),
	.Q(n_2345));
   AOI221_X2_50_SVT g78875__4319 (.A0(DPATH_RF_MEMORY_25__21_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__21_),
	.B1(FE_OFN53_n_1409),
	.C0(n_2275),
	.Q(n_2344));
   AOI221_X1_50_SVT g78876__8428 (.A0(DPATH_RF_MEMORY_28__16_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__16_),
	.B1(FE_OFN31_n_1379),
	.C0(n_2276),
	.Q(n_2343));
   NAND4T_X0_50_SVT g78877__5526 (.A(n_1492),
	.B(n_1491),
	.C(n_1495),
	.D(n_1493),
	.Q(n_2342));
   AOI221_X1_50_SVT g78878__6783 (.A0(DPATH_RF_MEMORY_9__10_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__10_),
	.B1(n_1417),
	.C0(n_2273),
	.Q(n_2341));
   AOI221_X1_50_SVT g78879__3680 (.A0(DPATH_RF_MEMORY_8__15_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__15_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2274),
	.Q(n_2340));
   NAND4_X2_50_SVT g78880__1617 (.A(n_1471),
	.B(n_1469),
	.C(n_2198),
	.D(n_2200),
	.Q(n_2339));
   NAND3T_X1_50_SVT g78881__2802 (.A(n_1990),
	.B(n_1988),
	.C(n_1992),
	.Q(n_2338));
   NAND3T_X0_50_SVT g78882__1705 (.A(n_2173),
	.B(n_2172),
	.C(n_2171),
	.Q(n_2337));
   NAND3T_X0_50_SVT g78883__5122 (.A(n_2154),
	.B(n_2153),
	.C(n_2152),
	.Q(n_2336));
   NAND3T_X1_50_SVT g78884__8246 (.A(n_2149),
	.B(n_2148),
	.C(n_2150),
	.Q(n_2335));
   NAND3_X2_50_SVT g78885__7098 (.A(n_2121),
	.B(n_2088),
	.C(n_2082),
	.Q(n_2334));
   NAND3T_X1_50_SVT g78886__6131 (.A(n_2130),
	.B(n_2132),
	.C(n_2134),
	.Q(n_2333));
   NAND3T_X1_50_SVT g78887__1881 (.A(n_2116),
	.B(n_2115),
	.C(n_2118),
	.Q(n_2332));
   NAND3T_X1_50_SVT g78888__5115 (.A(n_2113),
	.B(n_2111),
	.C(n_2114),
	.Q(n_2331));
   NAND3T_X1_50_SVT g78889__7482 (.A(n_2101),
	.B(n_2102),
	.C(n_2100),
	.Q(n_2330));
   NAND3_X2_50_SVT g78890__4733 (.A(n_2077),
	.B(n_2087),
	.C(n_2069),
	.Q(n_2329));
   NAND3T_X0_50_SVT g78891__6161 (.A(n_2083),
	.B(n_2086),
	.C(n_2084),
	.Q(n_2328));
   NAND3_X2_50_SVT g78892__9315 (.A(n_2120),
	.B(n_2109),
	.C(n_2095),
	.Q(n_2327));
   NAND3T_X1_50_SVT g78893__9945 (.A(n_2064),
	.B(n_2066),
	.C(n_2067),
	.Q(n_2326));
   NAND3_X2_50_SVT g78894__2883 (.A(n_2059),
	.B(n_2042),
	.C(n_2049),
	.Q(n_2325));
   NAND3_X2_50_SVT g78895__2346 (.A(n_2044),
	.B(n_2046),
	.C(n_2039),
	.Q(n_2324));
   NAND3T_X1_50_SVT g78896__1666 (.A(n_2045),
	.B(n_2043),
	.C(n_2047),
	.Q(n_2323));
   NAND3T_X1_50_SVT g78897__7410 (.A(n_2023),
	.B(n_2022),
	.C(n_2024),
	.Q(n_2322));
   NAND3_X2_50_SVT g78898__6417 (.A(n_2012),
	.B(n_1981),
	.C(n_1998),
	.Q(n_2321));
   NAND3T_X1_50_SVT g78899__5477 (.A(n_2005),
	.B(n_2004),
	.C(n_2007),
	.Q(n_2320));
   NAND3_X2_50_SVT g78900__2398 (.A(n_1993),
	.B(n_1987),
	.C(n_1989),
	.Q(n_2319));
   NAND3T_X1_50_SVT g78901__5107 (.A(n_2195),
	.B(n_2194),
	.C(n_2196),
	.Q(n_2318));
   NAND3T_X1_50_SVT g78902__6260 (.A(n_1968),
	.B(n_1967),
	.C(n_1969),
	.Q(n_2317));
   NAND3T_X1_50_SVT g78903__4319 (.A(n_1953),
	.B(n_1952),
	.C(n_2188),
	.Q(n_2316));
   NAND3_X2_50_SVT g78904__8428 (.A(n_1955),
	.B(n_1939),
	.C(n_1948),
	.Q(n_2315));
   NAND3T_X0_50_SVT g78905__5526 (.A(n_1944),
	.B(n_1942),
	.C(n_1941),
	.Q(n_2314));
   NAND3_X2_50_SVT g78906__6783 (.A(n_1927),
	.B(n_1630),
	.C(n_1925),
	.Q(n_2313));
   NAND3_X2_50_SVT g78907__3680 (.A(n_1913),
	.B(n_1911),
	.C(n_1908),
	.Q(n_2312));
   NAND3_X2_50_SVT g78908__1617 (.A(n_1905),
	.B(n_1903),
	.C(n_1902),
	.Q(n_2311));
   NAND3_X2_50_SVT g78909__2802 (.A(n_1896),
	.B(n_1893),
	.C(n_1890),
	.Q(n_2310));
   NAND3_X2_50_SVT g78910__1705 (.A(n_1892),
	.B(n_1891),
	.C(n_1889),
	.Q(n_2309));
   NAND3_X2_50_SVT g78911__5122 (.A(n_1880),
	.B(n_1872),
	.C(n_1864),
	.Q(n_2308));
   NAND3_X2_50_SVT g78912__8246 (.A(n_1868),
	.B(n_1867),
	.C(n_1866),
	.Q(n_2307));
   NAND3_X2_50_SVT g78913__7098 (.A(n_1833),
	.B(n_1801),
	.C(n_1805),
	.Q(n_2306));
   NAND3_X2_50_SVT g78914__6131 (.A(n_1850),
	.B(n_1843),
	.C(n_1848),
	.Q(n_2305));
   NAND3T_X1_50_SVT g78915__1881 (.A(n_1817),
	.B(n_1738),
	.C(n_1691),
	.Q(n_2304));
   NAND3_X2_50_SVT g78916__5115 (.A(n_1822),
	.B(n_1826),
	.C(n_1816),
	.Q(n_2303));
   NAND3_X2_50_SVT g78917__7482 (.A(n_1821),
	.B(n_1819),
	.C(n_1818),
	.Q(n_2302));
   NAND3T_X1_50_SVT g78918__4733 (.A(n_1770),
	.B(n_1771),
	.C(n_1775),
	.Q(n_2301));
   NAND3_X2_50_SVT g78919__6161 (.A(n_1772),
	.B(n_1768),
	.C(n_1764),
	.Q(n_2300));
   NAND3T_X1_50_SVT g78920__9315 (.A(n_1753),
	.B(n_1752),
	.C(n_1754),
	.Q(n_2299));
   NAND3T_X1_50_SVT g78921__9945 (.A(n_1729),
	.B(n_1730),
	.C(n_1728),
	.Q(n_2298));
   NAND3T_X1_50_SVT g78922__2883 (.A(n_1724),
	.B(n_1723),
	.C(n_1726),
	.Q(n_2297));
   NAND3T_X0_50_SVT g78923__2346 (.A(n_1713),
	.B(n_1715),
	.C(n_1714),
	.Q(n_2296));
   NAND3T_X1_50_SVT g78924__1666 (.A(n_1707),
	.B(n_1709),
	.C(n_1710),
	.Q(n_2295));
   NAND3_X2_50_SVT g78925__7410 (.A(n_1701),
	.B(n_1692),
	.C(n_1683),
	.Q(n_2294));
   NAND3T_X1_50_SVT g78926__6417 (.A(n_1697),
	.B(n_1694),
	.C(n_1698),
	.Q(n_2293));
   NAND3T_X1_50_SVT g78927__5477 (.A(n_1673),
	.B(n_1676),
	.C(n_1672),
	.Q(n_2292));
   NAND3_X2_50_SVT g78928__2398 (.A(n_1674),
	.B(n_1666),
	.C(n_1658),
	.Q(n_2291));
   NAND3_X2_50_SVT g78929__5107 (.A(n_1662),
	.B(n_1660),
	.C(n_1657),
	.Q(n_2290));
   NAND3T_X1_50_SVT g78930__6260 (.A(n_1650),
	.B(n_1786),
	.C(n_1652),
	.Q(n_2289));
   NAND3T_X1_50_SVT g78931__4319 (.A(n_1641),
	.B(n_1639),
	.C(n_1642),
	.Q(n_2288));
   NAND3T_X1_50_SVT g78932__8428 (.A(n_1618),
	.B(n_1863),
	.C(n_1620),
	.Q(n_2287));
   NAND3_X2_50_SVT g78933__5526 (.A(n_1609),
	.B(n_1598),
	.C(n_1596),
	.Q(n_2286));
   NAND3_X2_50_SVT g78934__6783 (.A(n_1601),
	.B(n_1589),
	.C(n_1595),
	.Q(n_2285));
   NAND3T_X1_50_SVT g78935__3680 (.A(n_1600),
	.B(n_1599),
	.C(n_1602),
	.Q(n_2284));
   NAND3T_X0_50_SVT g78936__1617 (.A(n_1580),
	.B(n_1578),
	.C(n_1577),
	.Q(n_2283));
   NAND3T_X1_50_SVT g78937__2802 (.A(n_1574),
	.B(n_1573),
	.C(n_1575),
	.Q(n_2282));
   NAND3T_X0_50_SVT g78938__1705 (.A(n_1563),
	.B(n_1562),
	.C(n_1561),
	.Q(n_2281));
   NAND3T_X1_50_SVT g78939__5122 (.A(n_1556),
	.B(n_1557),
	.C(n_1559),
	.Q(n_2280));
   NAND3T_X1_50_SVT g78940__8246 (.A(n_1542),
	.B(n_2065),
	.C(n_1543),
	.Q(n_2279));
   NAND3T_X1_50_SVT g78941__7098 (.A(n_2098),
	.B(n_1555),
	.C(n_2181),
	.Q(n_2278));
   NAND3T_X0_50_SVT g78942__6131 (.A(n_1527),
	.B(n_1526),
	.C(n_1525),
	.Q(n_2277));
   NAND3T_X0_50_SVT g78943__1881 (.A(n_1504),
	.B(n_1506),
	.C(n_1505),
	.Q(n_2276));
   NAND3_X2_50_SVT g78944__5115 (.A(n_1483),
	.B(n_1486),
	.C(n_1477),
	.Q(n_2275));
   NAND3T_X1_50_SVT g78945__7482 (.A(n_1487),
	.B(n_1485),
	.C(n_1488),
	.Q(n_2274));
   NAND3_X2_50_SVT g78946__4733 (.A(n_1484),
	.B(n_1472),
	.C(n_1479),
	.Q(n_2273));
   INV_A_OAI211_X2_50_SVT g78947__6161 (.A0(n_1394),
	.A1N(DPATH_RF_MEMORY_16__9_),
	.B0(n_2147),
	.C0(n_2145),
	.Q(n_2272));
   INV_A_OAI211_X2_50_SVT g78948__9315 (.A0(n_1394),
	.A1N(DPATH_RF_MEMORY_16__8_),
	.B0(n_2094),
	.C0(n_2091),
	.Q(n_2271));
   INV_A_OAI211_X2_50_SVT g78949__9945 (.A0(n_1428),
	.A1N(DPATH_RF_MEMORY_15__26_),
	.B0(n_2053),
	.C0(n_2040),
	.Q(n_2270));
   INV_A_OAI211_X2_50_SVT g78950__2883 (.A0(n_1426),
	.A1N(DPATH_RF_MEMORY_2__1_),
	.B0(n_1840),
	.C0(n_1839),
	.Q(n_2269));
   INV_A_OAI211_X2_50_SVT g78951__2346 (.A0(n_1373),
	.A1N(DPATH_RF_MEMORY_8__16_),
	.B0(n_1809),
	.C0(n_1811),
	.Q(n_2268));
   INV_A_OAI211_X2_50_SVT g78952__1666 (.A0(n_1332),
	.A1N(DPATH_RF_MEMORY_1__31_),
	.B0(n_1790),
	.C0(n_1789),
	.Q(n_2267));
   INV_A_OAI211_X2_50_SVT g78953__7410 (.A0(n_1426),
	.A1N(DPATH_RF_MEMORY_2__28_),
	.B0(n_1774),
	.C0(n_1781),
	.Q(n_2266));
   INV_A_OAI211_X2_50_SVT g78954__6417 (.A0(n_1373),
	.A1N(DPATH_RF_MEMORY_8__14_),
	.B0(n_1705),
	.C0(n_1708),
	.Q(n_2265));
   INV_A_OAI211_X2_50_SVT g78955__5477 (.A0(n_1416),
	.A1N(DPATH_RF_MEMORY_10__27_),
	.B0(n_1553),
	.C0(n_1541),
	.Q(n_2264));
   INV_A_OAI211_X2_50_SVT g78956__2398 (.A0(n_1373),
	.A1N(DPATH_RF_MEMORY_8__11_),
	.B0(n_1532),
	.C0(n_1536),
	.Q(n_2263));
   MUX2_X1_50_SVT g78957__5107 (.A(INSTR[9]),
	.B(INSTR[22]),
	.Q(DPATH_n_5228),
	.S0(n_2202));
   MUX2_X1_50_SVT g78958__6260 (.A(INSTR[10]),
	.B(INSTR[23]),
	.Q(DPATH_n_5227),
	.S0(n_2202));
   MUX2_X2_50_SVT g78959__4319 (.A(INSTR[11]),
	.B(INSTR[24]),
	.Q(DPATH_n_5226),
	.S0(n_2202));
   MUX2_X1_50_SVT g78960__8428 (.A(INSTR[8]),
	.B(INSTR[21]),
	.Q(DPATH_n_5229),
	.S0(n_2202));
   AOI221_X1_50_SVT g78962__6783 (.A0(DPATH_RF_MEMORY_9__26_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__26_),
	.B1(n_1399),
	.C0(n_1685),
	.Q(n_2262));
   AOI221_X1_50_SVT g78963__3680 (.A0(DPATH_RF_MEMORY_8__13_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__13_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2165),
	.Q(n_2261));
   AOI221_X1_50_SVT g78964__1617 (.A0(DPATH_RF_MEMORY_9__21_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__21_),
	.B1(n_1417),
	.C0(n_2163),
	.Q(n_2260));
   AOI221_X1_50_SVT g78965__2802 (.A0(DPATH_RF_MEMORY_13__11_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__11_),
	.B1(FE_OFN48_n_1401),
	.C0(n_2136),
	.Q(n_2259));
   AOI221_X1_50_SVT g78966__1705 (.A0(DPATH_RF_MEMORY_5__9_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__9_),
	.B1(FE_OFN49_n_1404),
	.C0(n_2096),
	.Q(n_2258));
   AOI221_X1_50_SVT g78967__5122 (.A0(DPATH_RF_MEMORY_12__8_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__8_),
	.B1(n_1450),
	.C0(n_2075),
	.Q(n_2257));
   AOI221_X1_50_SVT g78968__8246 (.A0(DPATH_RF_MEMORY_25__7_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__7_),
	.B1(FE_OFN38_n_1389),
	.C0(n_2055),
	.Q(n_2256));
   AOI221_X1_50_SVT g78969__7098 (.A0(DPATH_RF_MEMORY_25__6_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__6_),
	.B1(FE_OFN38_n_1389),
	.C0(n_2034),
	.Q(n_2255));
   AOI221_X0_50_SVT g78970__6131 (.A0(DPATH_RF_MEMORY_13__7_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__7_),
	.B1(n_1412),
	.C0(n_2018),
	.Q(n_2254));
   AOI221_X1_50_SVT g78971__1881 (.A0(DPATH_RF_MEMORY_4__5_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__5_),
	.B1(n_1446),
	.C0(n_2019),
	.Q(n_2253));
   AOI221_X1_50_SVT g78972__5115 (.A0(DPATH_RF_MEMORY_8__4_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__4_),
	.B1(FE_OFN69_n_1443),
	.C0(n_2000),
	.Q(n_2252));
   AOI221_X1_50_SVT g78973__7482 (.A0(DPATH_RF_MEMORY_12__3_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__3_),
	.B1(n_1450),
	.C0(n_2099),
	.Q(n_2251));
   AOI221_X0_50_SVT g78974__4733 (.A0(DPATH_RF_MEMORY_13__19_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__19_),
	.B1(n_1412),
	.C0(n_1963),
	.Q(n_2250));
   AOI221_X1_50_SVT g78975__6161 (.A0(DPATH_RF_MEMORY_25__2_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__2_),
	.B1(n_1389),
	.C0(n_2156),
	.Q(n_2249));
   AOI221_X0_50_SVT g78976__9315 (.A0(DPATH_RF_MEMORY_29__6_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__6_),
	.B1(FE_OFN29_n_1377),
	.C0(n_1965),
	.Q(n_2248));
   AOI221_X1_50_SVT g78977__9945 (.A0(DPATH_RF_MEMORY_25__1_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__1_),
	.B1(FE_OFN38_n_1389),
	.C0(n_1956),
	.Q(n_2247));
   AOI221_X1_50_SVT g78978__2883 (.A0(DPATH_RF_MEMORY_9__0_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__0_),
	.B1(n_1399),
	.C0(n_1932),
	.Q(n_2246));
   AOI221_X0_50_SVT g78979__2346 (.A0(DPATH_RF_MEMORY_13__5_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__5_),
	.B1(n_1412),
	.C0(n_1928),
	.Q(n_2245));
   AOI221_X1_50_SVT g78980__1666 (.A0(DPATH_RF_MEMORY_24__29_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__29_),
	.B1(FE_OFN33_n_1381),
	.C0(n_1920),
	.Q(n_2244));
   AOI221_X0_50_SVT g78981__7410 (.A0(DPATH_RF_MEMORY_24__18_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__18_),
	.B1(FE_OFN33_n_1381),
	.C0(n_1904),
	.Q(n_2243));
   AOI221_X0_50_SVT g78982__6417 (.A0(DPATH_RF_MEMORY_12__25_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__25_),
	.B1(FE_OFN40_n_1391),
	.C0(n_1894),
	.Q(n_2242));
   AOI221_X0_50_SVT g78983__5477 (.A0(DPATH_RF_MEMORY_25__3_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__3_),
	.B1(FE_OFN53_n_1409),
	.C0(n_1881),
	.Q(n_2241));
   AOI221_X0_50_SVT g78984__2398 (.A0(DPATH_RF_MEMORY_24__17_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__17_),
	.B1(FE_OFN33_n_1381),
	.C0(n_1857),
	.Q(n_2240));
   AOI221_X1_50_SVT g78985__5107 (.A0(DPATH_RF_MEMORY_29__2_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__2_),
	.B1(FE_OFN29_n_1377),
	.C0(n_1856),
	.Q(n_2239));
   AOI221_X1_50_SVT g78986__6260 (.A0(DPATH_RF_MEMORY_13__0_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__0_),
	.B1(n_1412),
	.C0(n_1828),
	.Q(n_2238));
   AOI221_X0_50_SVT g78987__4319 (.A0(DPATH_RF_MEMORY_12__15_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__15_),
	.B1(FE_OFN40_n_1391),
	.C0(n_1788),
	.Q(n_2237));
   AOI221_X0_50_SVT g78988__8428 (.A0(DPATH_RF_MEMORY_13__24_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__24_),
	.B1(n_1412),
	.C0(n_1773),
	.Q(n_2236));
   AOI221_X1_50_SVT g78989__5526 (.A0(DPATH_RF_MEMORY_29__30_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__30_),
	.B1(n_1378),
	.C0(n_1762),
	.Q(n_2235));
   AOI221_X1_50_SVT g78990__6783 (.A0(DPATH_RF_MEMORY_12__29_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__29_),
	.B1(n_1450),
	.C0(n_1742),
	.Q(n_2234));
   AOI221_X1_50_SVT g78991__3680 (.A0(DPATH_RF_MEMORY_12__14_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__14_),
	.B1(n_1450),
	.C0(n_2185),
	.Q(n_2233));
   AOI221_X1_50_SVT g78992__1617 (.A0(DPATH_RF_MEMORY_5__25_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__25_),
	.B1(FE_OFN49_n_1404),
	.C0(n_1668),
	.Q(n_2232));
   AOI221_X1_50_SVT g78993__2802 (.A0(DPATH_RF_MEMORY_12__24_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__24_),
	.B1(n_1450),
	.C0(n_1654),
	.Q(n_2231));
   AOI221_X0_50_SVT g78994__1705 (.A0(DPATH_RF_MEMORY_12__13_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__13_),
	.B1(FE_OFN40_n_1391),
	.C0(n_1631),
	.Q(n_2230));
   AOI221_X1_50_SVT g78995__5122 (.A0(DPATH_RF_MEMORY_28__23_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__23_),
	.B1(FE_OFN31_n_1379),
	.C0(n_1629),
	.Q(n_2229));
   AOI221_X0_50_SVT g78996__8246 (.A0(DPATH_RF_MEMORY_12__12_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__12_),
	.B1(FE_OFN40_n_1391),
	.C0(n_1616),
	.Q(n_2228));
   AOI221_X1_50_SVT g78997__7098 (.A0(DPATH_RF_MEMORY_13__22_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__22_),
	.B1(FE_OFN48_n_1401),
	.C0(n_1610),
	.Q(n_2227));
   AOI221_X1_50_SVT g78998__6131 (.A0(DPATH_RF_MEMORY_12__21_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__21_),
	.B1(n_1450),
	.C0(n_1590),
	.Q(n_2226));
   AOI221_X1_50_SVT g78999__1881 (.A0(DPATH_RF_MEMORY_24__30_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__30_),
	.B1(FE_OFN33_n_1381),
	.C0(n_1617),
	.Q(n_2225));
   AOI221_X1_50_SVT g79000__5115 (.A0(DPATH_RF_MEMORY_29__22_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__22_),
	.B1(FE_OFN29_n_1377),
	.C0(n_1544),
	.Q(n_2224));
   AOI221_X1_50_SVT g79001__7482 (.A0(DPATH_RF_MEMORY_4__18_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__18_),
	.B1(n_1446),
	.C0(n_1537),
	.Q(n_2223));
   AOI221_X1_50_SVT g79002__4733 (.A0(DPATH_RF_MEMORY_12__17_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__17_),
	.B1(n_1450),
	.C0(n_1517),
	.Q(n_2222));
   AOI221_X0_50_SVT g79003__6161 (.A0(DPATH_RF_MEMORY_4__10_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__10_),
	.B1(n_1420),
	.C0(n_1500),
	.Q(n_2221));
   AOI221_X1_50_SVT g79004__9315 (.A0(DPATH_RF_MEMORY_13__16_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__16_),
	.B1(FE_OFN48_n_1401),
	.C0(n_1497),
	.Q(n_2220));
   AOI221_X1_50_SVT g79005__9945 (.A0(DPATH_RF_MEMORY_29__15_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__15_),
	.B1(n_1378),
	.C0(n_1473),
	.Q(n_2219));
   AOI222_X1_50_SVT g79007__2346 (.A0(DPATH_RF_MEMORY_20__13_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_21__13_),
	.B1(n_1436),
	.C0(DPATH_RF_MEMORY_22__13_),
	.C1(n_1438),
	.Q(n_2218));
   AOI222_X1_50_SVT g79008__1666 (.A0(DPATH_RF_MEMORY_20__11_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_21__11_),
	.B1(FE_OFN64_n_1436),
	.C0(DPATH_RF_MEMORY_22__11_),
	.C1(FE_OFN65_n_1438),
	.Q(n_2217));
   AOI222_X1_50_SVT g79009__7410 (.A0(DPATH_RF_MEMORY_17__9_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_20__9_),
	.B1(n_1408),
	.C0(DPATH_RF_MEMORY_19__9_),
	.C1(n_1440),
	.Q(n_2216));
   AOI222_X1_50_SVT g79010__6417 (.A0(DPATH_RF_MEMORY_17__5_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_20__5_),
	.B1(n_1408),
	.C0(DPATH_RF_MEMORY_19__5_),
	.C1(n_1440),
	.Q(n_2215));
   AOI222_X1_50_SVT g79011__5477 (.A0(DPATH_RF_MEMORY_21__19_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__19_),
	.B1(FE_OFN25_n_1331),
	.C0(DPATH_RF_MEMORY_19__19_),
	.C1(FE_OFN44_n_1396),
	.Q(n_2214));
   AOI222_X1_50_SVT g79012__2398 (.A0(DPATH_RF_MEMORY_17__4_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_21__4_),
	.B1(FE_OFN64_n_1436),
	.C0(DPATH_RF_MEMORY_22__4_),
	.C1(FE_OFN65_n_1438),
	.Q(n_2213));
   AOI222_X1_50_SVT g79013__5107 (.A0(DPATH_RF_MEMORY_31__2_),
	.A1(n_1386),
	.B0(DPATH_RF_MEMORY_21__2_),
	.B1(n_1436),
	.C0(DPATH_RF_MEMORY_22__2_),
	.C1(FE_OFN65_n_1438),
	.Q(n_2212));
   AOI222_X1_50_SVT g79014__6260 (.A0(DPATH_RF_MEMORY_20__1_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_21__1_),
	.B1(n_1436),
	.C0(DPATH_RF_MEMORY_22__1_),
	.C1(FE_OFN65_n_1438),
	.Q(n_2211));
   AOI222_X1_50_SVT g79015__4319 (.A0(DPATH_RF_MEMORY_21__5_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__5_),
	.B1(FE_OFN25_n_1331),
	.C0(DPATH_RF_MEMORY_31__5_),
	.C1(FE_OFN35_n_1385),
	.Q(n_2210));
   AOI222_X1_50_SVT g79016__8428 (.A0(DPATH_RF_MEMORY_21__25_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__25_),
	.B1(FE_OFN25_n_1331),
	.C0(DPATH_RF_MEMORY_31__25_),
	.C1(FE_OFN35_n_1385),
	.Q(n_2209));
   AOI222_X1_50_SVT g79018__6783 (.A0(DPATH_RF_MEMORY_31__17_),
	.A1(FE_OFN35_n_1385),
	.B0(DPATH_RF_MEMORY_20__17_),
	.B1(FE_OFN41_n_1392),
	.C0(DPATH_RF_MEMORY_19__17_),
	.C1(FE_OFN44_n_1396),
	.Q(n_2207));
   AOI222_X1_50_SVT g79019__3680 (.A0(DPATH_RF_MEMORY_31__25_),
	.A1(FE_OFN36_n_1386),
	.B0(DPATH_RF_MEMORY_21__25_),
	.B1(FE_OFN64_n_1436),
	.C0(DPATH_RF_MEMORY_22__25_),
	.C1(FE_OFN65_n_1438),
	.Q(n_2206));
   AOI222_X1_50_SVT g79020__1617 (.A0(DPATH_RF_MEMORY_17__24_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_20__24_),
	.B1(FE_OFN52_n_1408),
	.C0(DPATH_RF_MEMORY_19__24_),
	.C1(FE_OFN66_n_1440),
	.Q(n_2205));
   AOI222_X1_50_SVT g79021__2802 (.A0(DPATH_RF_MEMORY_21__18_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__18_),
	.B1(FE_OFN65_n_1438),
	.C0(DPATH_RF_MEMORY_19__18_),
	.C1(FE_OFN66_n_1440),
	.Q(n_2204));
   AOI222_X1_50_SVT g79022__1705 (.A0(DPATH_RF_MEMORY_22__18_),
	.A1(FE_OFN25_n_1331),
	.B0(DPATH_RF_MEMORY_20__18_),
	.B1(FE_OFN41_n_1392),
	.C0(DPATH_RF_MEMORY_19__18_),
	.C1(FE_OFN44_n_1396),
	.Q(n_2203));
   AOI22_X1_50_SVT g79023__5122 (.A0(DPATH_RF_MEMORY_20__16_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__16_),
	.B1(FE_OFN44_n_1396),
	.Q(n_2201));
   AOI22_X1_50_SVT g79024__8246 (.A0(DPATH_RF_MEMORY_8__14_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__14_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2200));
   AOI22_X1_50_SVT g79025__7098 (.A0(DPATH_RF_MEMORY_21__21_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__21_),
	.B1(FE_OFN25_n_1331),
	.Q(n_2199));
   AOI22_X1_50_SVT g79026__6131 (.A0(DPATH_RF_MEMORY_1__14_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__14_),
	.B1(n_1434),
	.Q(n_2198));
   AOI22_X1_50_SVT g79027__1881 (.A0(DPATH_RF_MEMORY_29__10_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__10_),
	.B1(n_1377),
	.Q(n_2197));
   AOI22_X1_50_SVT g79028__5115 (.A0(DPATH_RF_MEMORY_24__14_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__14_),
	.B1(n_1445),
	.Q(n_2196));
   AOI22_X1_50_SVT g79029__7482 (.A0(DPATH_RF_MEMORY_28__14_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__14_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2195));
   AOI22_X1_50_SVT g79030__4733 (.A0(DPATH_RF_MEMORY_25__14_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__14_),
	.B1(FE_OFN38_n_1389),
	.Q(n_2194));
   AOI22_X1_50_SVT g79031__6161 (.A0(DPATH_RF_MEMORY_17__26_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__26_),
	.B1(FE_OFN57_n_1419),
	.Q(n_2193));
   AOI22_X1_50_SVT g79032__9315 (.A0(DPATH_RF_MEMORY_28__10_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__10_),
	.B1(FE_OFN55_n_1413),
	.Q(n_2192));
   AOI22_X1_50_SVT g79033__9945 (.A0(DPATH_RF_MEMORY_17__14_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__14_),
	.B1(FE_OFN36_n_1386),
	.Q(n_2191));
   AOI22_X1_50_SVT g79034__2883 (.A0(DPATH_RF_MEMORY_25__10_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__10_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2190));
   AOI22_X1_50_SVT g79035__2346 (.A0(DPATH_RF_MEMORY_21__14_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__14_),
	.B1(FE_OFN65_n_1438),
	.Q(n_2189));
   AOI22_X1_50_SVT g79036__1666 (.A0(DPATH_RF_MEMORY_4__1_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__1_),
	.B1(n_1446),
	.Q(n_2188));
   AOI22_X1_50_SVT g79037__7410 (.A0(DPATH_RF_MEMORY_16__14_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__14_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2187));
   AOI22_X1_50_SVT g79038__6417 (.A0(DPATH_RF_MEMORY_9__14_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__14_),
	.B1(n_1399),
	.Q(n_2186));
   AO22_X0_50_SVT g79039__5477 (.A0(DPATH_RF_MEMORY_13__14_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__14_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2185));
   AOI22_X1_50_SVT g79040__2398 (.A0(DPATH_RF_MEMORY_24__10_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__10_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2184));
   AOI22_X1_50_SVT g79041__5107 (.A0(DPATH_RF_MEMORY_17__21_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__21_),
	.B1(FE_OFN35_n_1385),
	.Q(n_2183));
   AOI22_X1_50_SVT g79042__6260 (.A0(DPATH_RF_MEMORY_17__13_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_19__13_),
	.B1(n_1440),
	.Q(n_2182));
   AOI22_X1_50_SVT g79043__4319 (.A0(DPATH_RF_MEMORY_5__31_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__31_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2181));
   AOI22_X1_50_SVT g79044__8428 (.A0(DPATH_RF_MEMORY_17__9_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_18__9_),
	.B1(FE_OFN57_n_1419),
	.Q(n_2180));
   AOI22_X1_50_SVT g79045__5526 (.A0(DPATH_RF_MEMORY_9__13_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__13_),
	.B1(n_1399),
	.Q(n_2179));
   AOI22_X1_50_SVT g79046__6783 (.A0(DPATH_RF_MEMORY_12__13_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__13_),
	.B1(n_1450),
	.Q(n_2178));
   AOI22_X1_50_SVT g79047__3680 (.A0(DPATH_RF_MEMORY_13__21_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__21_),
	.B1(n_1412),
	.Q(n_2177));
   AOI22_X1_50_SVT g79048__1617 (.A0(DPATH_RF_MEMORY_13__13_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__13_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2176));
   AOI22_X1_50_SVT g79049__2802 (.A0(DPATH_RF_MEMORY_16__13_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__13_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2175));
   AOI22_X1_50_SVT g79050__1705 (.A0(DPATH_RF_MEMORY_20__9_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__9_),
	.B1(FE_OFN44_n_1396),
	.Q(n_2174));
   AOI22_X1_50_SVT g79051__5122 (.A0(DPATH_RF_MEMORY_25__13_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__13_),
	.B1(n_1389),
	.Q(n_2173));
   AOI22_X1_50_SVT g79052__8246 (.A0(DPATH_RF_MEMORY_29__13_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__13_),
	.B1(n_1378),
	.Q(n_2172));
   AOI22_X1_50_SVT g79053__7098 (.A0(DPATH_RF_MEMORY_28__13_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__13_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2171));
   AO22_X0_50_SVT g79054__6131 (.A0(DPATH_RF_MEMORY_20__26_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__26_),
	.B1(FE_OFN44_n_1396),
	.Q(n_2170));
   AOI22_X1_50_SVT g79055__1881 (.A0(DPATH_RF_MEMORY_5__13_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__13_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2169));
   AOI22_X1_50_SVT g79056__5115 (.A0(DPATH_RF_MEMORY_12__21_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__21_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2168));
   AOI22_X1_50_SVT g79057__7482 (.A0(DPATH_RF_MEMORY_1__13_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__13_),
	.B1(n_1434),
	.Q(n_2167));
   AOI22_X1_50_SVT g79058__4733 (.A0(DPATH_RF_MEMORY_24__9_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__9_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2166));
   AO22_X0_50_SVT g79059__6161 (.A0(DPATH_RF_MEMORY_4__13_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__13_),
	.B1(n_1446),
	.Q(n_2165));
   AO22_X0_50_SVT g79060__9315 (.A0(DPATH_RF_MEMORY_22__12_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_19__12_),
	.B1(FE_OFN66_n_1440),
	.Q(n_2164));
   AO22_X0_50_SVT g79061__9945 (.A0(DPATH_RF_MEMORY_16__21_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__21_),
	.B1(FE_OFN62_n_1429),
	.Q(n_2163));
   AOI22_X1_50_SVT g79062__2883 (.A0(DPATH_RF_MEMORY_28__12_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__12_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2162));
   AOI22_X1_50_SVT g79063__2346 (.A0(DPATH_RF_MEMORY_28__9_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__9_),
	.B1(FE_OFN55_n_1413),
	.Q(n_2161));
   AOI22_X1_50_SVT g79064__1666 (.A0(DPATH_RF_MEMORY_29__12_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__12_),
	.B1(n_1378),
	.Q(n_2160));
   AOI22_X1_50_SVT g79065__7410 (.A0(DPATH_RF_MEMORY_29__9_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__9_),
	.B1(FE_OFN29_n_1377),
	.Q(n_2159));
   AOI22_X1_50_SVT g79066__6417 (.A0(DPATH_RF_MEMORY_25__12_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__12_),
	.B1(FE_OFN38_n_1389),
	.Q(n_2158));
   AOI22_X1_50_SVT g79067__5477 (.A0(DPATH_RF_MEMORY_24__12_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__12_),
	.B1(n_1445),
	.Q(n_2157));
   AO22_X0_50_SVT g79068__2398 (.A0(DPATH_RF_MEMORY_28__2_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__2_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2156));
   AOI22_X1_50_SVT g79069__5107 (.A0(DPATH_RF_MEMORY_25__9_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__9_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2155));
   AOI22_X1_50_SVT g79070__6260 (.A0(DPATH_RF_MEMORY_12__12_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__12_),
	.B1(n_1450),
	.Q(n_2154));
   AOI22_X1_50_SVT g79071__4319 (.A0(DPATH_RF_MEMORY_13__12_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__12_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2153));
   AOI22_X1_50_SVT g79072__8428 (.A0(DPATH_RF_MEMORY_16__12_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__12_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2152));
   AOI22_X1_50_SVT g79073__5526 (.A0(DPATH_RF_MEMORY_21__26_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__26_),
	.B1(FE_OFN25_n_1331),
	.Q(n_2151));
   AOI22_X1_50_SVT g79074__6783 (.A0(DPATH_RF_MEMORY_1__12_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__12_),
	.B1(n_1434),
	.Q(n_2150));
   AOI22_X1_50_SVT g79075__3680 (.A0(DPATH_RF_MEMORY_5__12_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__12_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2149));
   AOI22_X1_50_SVT g79076__1617 (.A0(DPATH_RF_MEMORY_8__12_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__12_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2148));
   AOI22_X1_50_SVT g79077__2802 (.A0(DPATH_RF_MEMORY_13__9_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__9_),
	.B1(n_1412),
	.Q(n_2147));
   AOI22_X1_50_SVT g79078__1705 (.A0(DPATH_RF_MEMORY_17__11_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_19__11_),
	.B1(FE_OFN66_n_1440),
	.Q(n_2146));
   AOI22_X1_50_SVT g79079__5122 (.A0(DPATH_RF_MEMORY_9__9_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__9_),
	.B1(n_1417),
	.Q(n_2145));
   AOI22_X1_50_SVT g79080__8246 (.A0(DPATH_RF_MEMORY_28__11_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__11_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2144));
   AOI22_X1_50_SVT g79081__7098 (.A0(DPATH_RF_MEMORY_29__11_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__11_),
	.B1(n_1378),
	.Q(n_2143));
   AOI22_X1_50_SVT g79082__6131 (.A0(DPATH_RF_MEMORY_8__9_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__9_),
	.B1(n_1403),
	.Q(n_2142));
   AOI22_X1_50_SVT g79083__1881 (.A0(DPATH_RF_MEMORY_25__11_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__11_),
	.B1(FE_OFN38_n_1389),
	.Q(n_2141));
   AOI22_X1_50_SVT g79084__5115 (.A0(DPATH_RF_MEMORY_24__11_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__11_),
	.B1(n_1445),
	.Q(n_2140));
   AOI22_X1_50_SVT g79085__7482 (.A0(DPATH_RF_MEMORY_9__11_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__11_),
	.B1(n_1399),
	.Q(n_2139));
   AOI22_X1_50_SVT g79086__4733 (.A0(DPATH_RF_MEMORY_13__20_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__20_),
	.B1(n_1412),
	.Q(n_2138));
   AOI22_X1_50_SVT g79087__6161 (.A0(DPATH_RF_MEMORY_1__9_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__9_),
	.B1(n_1427),
	.Q(n_2137));
   AO22_X0_50_SVT g79088__9315 (.A0(DPATH_RF_MEMORY_16__11_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__11_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2136));
   AOI22_X1_50_SVT g79089__9945 (.A0(DPATH_RF_MEMORY_5__9_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__9_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2135));
   AOI22_X1_50_SVT g79090__2883 (.A0(DPATH_RF_MEMORY_5__11_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__11_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2134));
   AOI22_X1_50_SVT g79091__2346 (.A0(DPATH_RF_MEMORY_12__20_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__20_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2133));
   AOI22_X1_50_SVT g79092__1666 (.A0(DPATH_RF_MEMORY_8__11_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__11_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2132));
   AOI22_X1_50_SVT g79093__7410 (.A0(DPATH_RF_MEMORY_4__9_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__9_),
	.B1(n_1420),
	.Q(n_2131));
   AOI22_X1_50_SVT g79094__6417 (.A0(DPATH_RF_MEMORY_4__11_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__11_),
	.B1(n_1446),
	.Q(n_2130));
   AOI22_X1_50_SVT g79095__5477 (.A0(DPATH_RF_MEMORY_13__18_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__18_),
	.B1(n_1412),
	.Q(n_2129));
   AOI22_X1_50_SVT g79096__2398 (.A0(DPATH_RF_MEMORY_13__10_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__10_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2128));
   AOI22_X1_50_SVT g79097__5107 (.A0(DPATH_RF_MEMORY_17__8_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_18__8_),
	.B1(FE_OFN57_n_1419),
	.Q(n_2127));
   AOI22_X1_50_SVT g79098__6260 (.A0(DPATH_RF_MEMORY_12__10_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__10_),
	.B1(n_1450),
	.Q(n_2126));
   AOI22_X1_50_SVT g79099__4319 (.A0(DPATH_RF_MEMORY_16__10_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__10_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2125));
   AOI22_X1_50_SVT g79100__8428 (.A0(DPATH_RF_MEMORY_9__10_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__10_),
	.B1(n_1399),
	.Q(n_2124));
   AOI22_X1_50_SVT g79101__5526 (.A0(DPATH_RF_MEMORY_25__29_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__29_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2123));
   AOI22_X1_50_SVT g79102__6783 (.A0(DPATH_RF_MEMORY_16__20_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__20_),
	.B1(FE_OFN62_n_1429),
	.Q(n_2122));
   AOI22_X1_50_SVT g79103__3680 (.A0(DPATH_RF_MEMORY_1__29_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__29_),
	.B1(n_1427),
	.Q(n_2121));
   AOI22_X1_50_SVT g79104__1617 (.A0(DPATH_RF_MEMORY_29__26_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__26_),
	.B1(FE_OFN29_n_1377),
	.Q(n_2120));
   AOI22_X1_50_SVT g79105__2802 (.A0(DPATH_RF_MEMORY_20__8_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__8_),
	.B1(FE_OFN44_n_1396),
	.Q(n_2119));
   AOI22_X1_50_SVT g79106__1705 (.A0(DPATH_RF_MEMORY_24__10_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__10_),
	.B1(n_1445),
	.Q(n_2118));
   AOI22_X1_50_SVT g79107__5122 (.A0(DPATH_RF_MEMORY_9__20_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__20_),
	.B1(n_1417),
	.Q(n_2117));
   AOI22_X1_50_SVT g79108__8246 (.A0(DPATH_RF_MEMORY_28__10_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__10_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2116));
   AOI22_X1_50_SVT g79109__7098 (.A0(DPATH_RF_MEMORY_25__10_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__10_),
	.B1(n_1389),
	.Q(n_2115));
   AOI22_X1_50_SVT g79110__6131 (.A0(DPATH_RF_MEMORY_1__10_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__10_),
	.B1(n_1434),
	.Q(n_2114));
   AOI22_X1_50_SVT g79111__1881 (.A0(DPATH_RF_MEMORY_5__10_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__10_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2113));
   AOI22_X1_50_SVT g79112__5115 (.A0(DPATH_RF_MEMORY_28__8_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__8_),
	.B1(FE_OFN55_n_1413),
	.Q(n_2112));
   AOI22_X1_50_SVT g79113__7482 (.A0(DPATH_RF_MEMORY_4__10_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__10_),
	.B1(n_1446),
	.Q(n_2111));
   AOI22_X1_50_SVT g79114__4733 (.A0(DPATH_RF_MEMORY_22__9_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_31__9_),
	.B1(n_1386),
	.Q(n_2110));
   AOI22_X1_50_SVT g79115__6161 (.A0(DPATH_RF_MEMORY_25__26_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__26_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2109));
   AOI22_X1_50_SVT g79116__9315 (.A0(DPATH_RF_MEMORY_29__8_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__8_),
	.B1(FE_OFN29_n_1377),
	.Q(n_2108));
   AOI22_X1_50_SVT g79117__9945 (.A0(DPATH_RF_MEMORY_24__9_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__9_),
	.B1(n_1445),
	.Q(n_2107));
   AOI22_X1_50_SVT g79118__2883 (.A0(DPATH_RF_MEMORY_25__9_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__9_),
	.B1(FE_OFN38_n_1389),
	.Q(n_2106));
   AOI22_X1_50_SVT g79119__2346 (.A0(DPATH_RF_MEMORY_25__8_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__8_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2105));
   AOI22_X1_50_SVT g79120__1666 (.A0(DPATH_RF_MEMORY_24__8_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__8_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2104));
   AOI22_X1_50_SVT g79121__7410 (.A0(DPATH_RF_MEMORY_28__9_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__9_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2103));
   AOI22_X1_50_SVT g79122__6417 (.A0(DPATH_RF_MEMORY_16__9_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__9_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2102));
   AOI22_X1_50_SVT g79123__5477 (.A0(DPATH_RF_MEMORY_12__9_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__9_),
	.B1(n_1450),
	.Q(n_2101));
   AOI22_X1_50_SVT g79124__2398 (.A0(DPATH_RF_MEMORY_9__9_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__9_),
	.B1(n_1399),
	.Q(n_2100));
   AO22_X0_50_SVT g79125__5107 (.A0(DPATH_RF_MEMORY_13__3_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__3_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2099));
   AOI22_X1_50_SVT g79126__6260 (.A0(DPATH_RF_MEMORY_1__31_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__31_),
	.B1(n_1427),
	.Q(n_2098));
   AOI22_X1_50_SVT g79127__4319 (.A0(DPATH_RF_MEMORY_8__9_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__9_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2097));
   AO22_X0_50_SVT g79128__8428 (.A0(DPATH_RF_MEMORY_1__9_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__9_),
	.B1(n_1434),
	.Q(n_2096));
   AOI22_X1_50_SVT g79129__5526 (.A0(DPATH_RF_MEMORY_24__26_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__26_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2095));
   AOI22_X1_50_SVT g79130__6783 (.A0(DPATH_RF_MEMORY_12__8_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__8_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2094));
   AOI22_X1_50_SVT g79131__3680 (.A0(DPATH_RF_MEMORY_8__8_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__8_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2093));
   AOI22_X1_50_SVT g79132__1617 (.A0(DPATH_RF_MEMORY_1__8_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__8_),
	.B1(n_1434),
	.Q(n_2092));
   AOI22_X1_50_SVT g79133__2802 (.A0(DPATH_RF_MEMORY_9__8_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__8_),
	.B1(n_1417),
	.Q(n_2091));
   AOI22_X1_50_SVT g79134__1705 (.A0(DPATH_RF_MEMORY_5__8_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__8_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2090));
   AOI22_X1_50_SVT g79135__5122 (.A0(DPATH_RF_MEMORY_4__8_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__8_),
	.B1(n_1446),
	.Q(n_2089));
   AOI22_X1_50_SVT g79136__8246 (.A0(DPATH_RF_MEMORY_5__29_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__29_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2088));
   AOI22_X1_50_SVT g79137__7098 (.A0(DPATH_RF_MEMORY_24__20_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__20_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2087));
   AOI22_X1_50_SVT g79138__6131 (.A0(DPATH_RF_MEMORY_29__8_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__8_),
	.B1(n_1378),
	.Q(n_2086));
   AOI22_X1_50_SVT g79139__1881 (.A0(DPATH_RF_MEMORY_4__8_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__8_),
	.B1(n_1420),
	.Q(n_2085));
   AOI22_X1_50_SVT g79140__5115 (.A0(DPATH_RF_MEMORY_28__8_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__8_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2084));
   AOI22_X1_50_SVT g79141__7482 (.A0(DPATH_RF_MEMORY_24__8_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__8_),
	.B1(n_1445),
	.Q(n_2083));
   AOI22_X1_50_SVT g79142__4733 (.A0(DPATH_RF_MEMORY_4__29_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__29_),
	.B1(n_1420),
	.Q(n_2082));
   AOI22_X1_50_SVT g79143__6161 (.A0(DPATH_RF_MEMORY_17__8_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__8_),
	.B1(n_1386),
	.Q(n_2081));
   AOI22_X1_50_SVT g79144__9315 (.A0(DPATH_RF_MEMORY_5__8_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__8_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2080));
   AOI22_X1_50_SVT g79145__9945 (.A0(DPATH_RF_MEMORY_21__8_),
	.A1(n_1436),
	.B0(DPATH_RF_MEMORY_22__8_),
	.B1(FE_OFN65_n_1438),
	.Q(n_2079));
   AOI22_X1_50_SVT g79146__2883 (.A0(DPATH_RF_MEMORY_16__8_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__8_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2078));
   AOI22_X1_50_SVT g79147__2346 (.A0(DPATH_RF_MEMORY_29__20_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__20_),
	.B1(FE_OFN29_n_1377),
	.Q(n_2077));
   AOI22_X1_50_SVT g79148__1666 (.A0(DPATH_RF_MEMORY_9__8_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__8_),
	.B1(n_1399),
	.Q(n_2076));
   AO22_X0_50_SVT g79149__7410 (.A0(DPATH_RF_MEMORY_13__8_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__8_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2075));
   AOI22_X1_50_SVT g79150__6417 (.A0(DPATH_RF_MEMORY_9__7_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__7_),
	.B1(n_1399),
	.Q(n_2074));
   AOI22_X1_50_SVT g79151__5477 (.A0(DPATH_RF_MEMORY_12__7_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__7_),
	.B1(n_1450),
	.Q(n_2073));
   AOI22_X1_50_SVT g79152__2398 (.A0(DPATH_RF_MEMORY_1__8_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__8_),
	.B1(n_1427),
	.Q(n_2072));
   AOI22_X1_50_SVT g79153__5107 (.A0(DPATH_RF_MEMORY_13__7_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__7_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2071));
   AOI22_X1_50_SVT g79154__6260 (.A0(DPATH_RF_MEMORY_16__7_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__7_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2070));
   AOI22_X1_50_SVT g79155__4319 (.A0(DPATH_RF_MEMORY_28__20_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__20_),
	.B1(FE_OFN55_n_1413),
	.Q(n_2069));
   AOI22_X1_50_SVT g79156__8428 (.A0(DPATH_RF_MEMORY_5__7_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__7_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2068));
   AOI22_X1_50_SVT g79157__5526 (.A0(DPATH_RF_MEMORY_5__7_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__7_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2067));
   AOI22_X1_50_SVT g79158__6783 (.A0(DPATH_RF_MEMORY_8__7_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__7_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2066));
   AOI22_X1_50_SVT g79159__3680 (.A0(DPATH_RF_MEMORY_25__18_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__18_),
	.B1(n_1389),
	.Q(n_2065));
   AOI22_X1_50_SVT g79160__1617 (.A0(DPATH_RF_MEMORY_4__7_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__7_),
	.B1(n_1446),
	.Q(n_2064));
   AOI22_X1_50_SVT g79161__2802 (.A0(DPATH_RF_MEMORY_21__7_),
	.A1(n_1436),
	.B0(DPATH_RF_MEMORY_22__7_),
	.B1(FE_OFN65_n_1438),
	.Q(n_2063));
   AOI22_X1_50_SVT g79162__1705 (.A0(DPATH_RF_MEMORY_1__7_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__7_),
	.B1(n_1427),
	.Q(n_2062));
   AOI22_X1_50_SVT g79163__5122 (.A0(DPATH_RF_MEMORY_8__7_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__7_),
	.B1(n_1403),
	.Q(n_2061));
   AOI22_X1_50_SVT g79164__8246 (.A0(DPATH_RF_MEMORY_17__7_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__7_),
	.B1(n_1386),
	.Q(n_2060));
   AOI22_X1_50_SVT g79165__7098 (.A0(DPATH_RF_MEMORY_4__20_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__20_),
	.B1(n_1420),
	.Q(n_2059));
   AOI22_X1_50_SVT g79166__6131 (.A0(DPATH_RF_MEMORY_24__7_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__7_),
	.B1(n_1445),
	.Q(n_2058));
   AOI22_X1_50_SVT g79167__1881 (.A0(DPATH_RF_MEMORY_4__7_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__7_),
	.B1(n_1420),
	.Q(n_2057));
   AOI22_X1_50_SVT g79168__5115 (.A0(DPATH_RF_MEMORY_29__7_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__7_),
	.B1(n_1378),
	.Q(n_2056));
   AO22_X0_50_SVT g79169__7482 (.A0(DPATH_RF_MEMORY_28__7_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__7_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2055));
   AOI22_X1_50_SVT g79170__4733 (.A0(DPATH_RF_MEMORY_22__5_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_31__5_),
	.B1(n_1386),
	.Q(n_2054));
   AOI22_X1_50_SVT g79171__6161 (.A0(DPATH_RF_MEMORY_12__26_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__26_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2053));
   AOI22_X1_50_SVT g79172__9315 (.A0(DPATH_RF_MEMORY_16__6_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__6_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2052));
   AOI22_X1_50_SVT g79173__9945 (.A0(DPATH_RF_MEMORY_9__6_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__6_),
	.B1(n_1399),
	.Q(n_2051));
   AOI22_X1_50_SVT g79174__2883 (.A0(DPATH_RF_MEMORY_13__6_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__6_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2050));
   AOI22_X1_50_SVT g79175__2346 (.A0(DPATH_RF_MEMORY_5__20_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__20_),
	.B1(FE_OFN59_n_1423),
	.Q(n_2049));
   AOI22_X1_50_SVT g79176__1666 (.A0(DPATH_RF_MEMORY_12__6_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__6_),
	.B1(n_1450),
	.Q(n_2048));
   AOI22_X1_50_SVT g79177__7410 (.A0(DPATH_RF_MEMORY_8__6_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__6_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2047));
   AOI22_X1_50_SVT g79178__6417 (.A0(DPATH_RF_MEMORY_28__7_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__7_),
	.B1(FE_OFN55_n_1413),
	.Q(n_2046));
   AOI22_X1_50_SVT g79179__5477 (.A0(DPATH_RF_MEMORY_5__6_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__6_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2045));
   AOI22_X1_50_SVT g79180__2398 (.A0(DPATH_RF_MEMORY_29__7_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__7_),
	.B1(FE_OFN29_n_1377),
	.Q(n_2044));
   AOI22_X1_50_SVT g79181__5107 (.A0(DPATH_RF_MEMORY_1__6_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__6_),
	.B1(n_1434),
	.Q(n_2043));
   AOI22_X1_50_SVT g79182__6260 (.A0(DPATH_RF_MEMORY_8__20_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__20_),
	.B1(n_1403),
	.Q(n_2042));
   AOI22_X1_50_SVT g79183__4319 (.A0(DPATH_RF_MEMORY_21__6_),
	.A1(n_1436),
	.B0(DPATH_RF_MEMORY_22__6_),
	.B1(FE_OFN65_n_1438),
	.Q(n_2041));
   AOI22_X1_50_SVT g79184__8428 (.A0(DPATH_RF_MEMORY_9__26_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__26_),
	.B1(n_1417),
	.Q(n_2040));
   AOI22_X1_50_SVT g79185__5526 (.A0(DPATH_RF_MEMORY_25__7_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__7_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2039));
   AOI22_X1_50_SVT g79186__6783 (.A0(DPATH_RF_MEMORY_20__6_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_19__6_),
	.B1(n_1440),
	.Q(n_2038));
   AOI22_X1_50_SVT g79187__3680 (.A0(DPATH_RF_MEMORY_29__6_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__6_),
	.B1(n_1378),
	.Q(n_2037));
   AOI22_X1_50_SVT g79188__1617 (.A0(DPATH_RF_MEMORY_21__7_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__7_),
	.B1(FE_OFN25_n_1331),
	.Q(n_2036));
   AOI22_X1_50_SVT g79189__2802 (.A0(DPATH_RF_MEMORY_24__6_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__6_),
	.B1(n_1445),
	.Q(n_2035));
   AO22_X0_50_SVT g79190__1705 (.A0(DPATH_RF_MEMORY_28__6_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__6_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2034));
   AOI22_X1_50_SVT g79191__5122 (.A0(DPATH_RF_MEMORY_20__19_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_31__19_),
	.B1(FE_OFN35_n_1385),
	.Q(n_2033));
   AOI22_X1_50_SVT g79192__8246 (.A0(DPATH_RF_MEMORY_20__29_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__29_),
	.B1(FE_OFN44_n_1396),
	.Q(n_2032));
   AOI22_X1_50_SVT g79193__7098 (.A0(DPATH_RF_MEMORY_18__7_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__7_),
	.B1(FE_OFN35_n_1385),
	.Q(n_2031));
   AOI22_X1_50_SVT g79194__6131 (.A0(DPATH_RF_MEMORY_9__5_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__5_),
	.B1(n_1399),
	.Q(n_2030));
   AOI22_X1_50_SVT g79195__1881 (.A0(DPATH_RF_MEMORY_16__5_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__5_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2029));
   AOI22_X1_50_SVT g79196__5115 (.A0(DPATH_RF_MEMORY_13__5_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__5_),
	.B1(FE_OFN48_n_1401),
	.Q(n_2028));
   AOI22_X1_50_SVT g79197__7482 (.A0(DPATH_RF_MEMORY_12__5_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__5_),
	.B1(n_1450),
	.Q(n_2027));
   AOI22_X1_50_SVT g79198__4733 (.A0(DPATH_RF_MEMORY_12__7_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__7_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2026));
   AOI22_X1_50_SVT g79199__6161 (.A0(DPATH_RF_MEMORY_9__7_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__7_),
	.B1(n_1417),
	.Q(n_2025));
   AOI22_X1_50_SVT g79200__9315 (.A0(DPATH_RF_MEMORY_25__5_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__5_),
	.B1(n_1389),
	.Q(n_2024));
   AOI22_X1_50_SVT g79201__9945 (.A0(DPATH_RF_MEMORY_28__5_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__5_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2023));
   AOI22_X1_50_SVT g79202__2883 (.A0(DPATH_RF_MEMORY_24__5_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__5_),
	.B1(n_1445),
	.Q(n_2022));
   AOI22_X1_50_SVT g79203__2346 (.A0(DPATH_RF_MEMORY_8__5_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__5_),
	.B1(FE_OFN69_n_1443),
	.Q(n_2021));
   AOI22_X1_50_SVT g79204__1666 (.A0(DPATH_RF_MEMORY_1__5_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__5_),
	.B1(n_1434),
	.Q(n_2020));
   AO22_X0_50_SVT g79205__7410 (.A0(DPATH_RF_MEMORY_5__5_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__5_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2019));
   AO22_X0_50_SVT g79206__6417 (.A0(DPATH_RF_MEMORY_16__7_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__7_),
	.B1(FE_OFN62_n_1429),
	.Q(n_2018));
   AOI22_X1_50_SVT g79207__5477 (.A0(DPATH_RF_MEMORY_20__4_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_31__4_),
	.B1(FE_OFN36_n_1386),
	.Q(n_2017));
   AOI22_X1_50_SVT g79208__2398 (.A0(DPATH_RF_MEMORY_16__3_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__3_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2016));
   AOI22_X1_50_SVT g79209__5107 (.A0(DPATH_RF_MEMORY_25__19_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__19_),
	.B1(FE_OFN53_n_1409),
	.Q(n_2015));
   AOI22_X1_50_SVT g79210__6260 (.A0(DPATH_RF_MEMORY_12__4_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__4_),
	.B1(n_1450),
	.Q(n_2014));
   AOI22_X1_50_SVT g79211__4319 (.A0(DPATH_RF_MEMORY_4__9_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__9_),
	.B1(n_1446),
	.Q(n_2013));
   AOI22_X1_50_SVT g79212__8428 (.A0(DPATH_RF_MEMORY_8__26_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__26_),
	.B1(n_1403),
	.Q(n_2012));
   AOI22_X1_50_SVT g79213__5526 (.A0(DPATH_RF_MEMORY_13__6_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__6_),
	.B1(n_1412),
	.Q(n_2011));
   AOI22_X1_50_SVT g79214__6783 (.A0(DPATH_RF_MEMORY_16__4_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__4_),
	.B1(FE_OFN72_n_1448),
	.Q(n_2010));
   AOI22_X1_50_SVT g79215__3680 (.A0(DPATH_RF_MEMORY_24__19_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__19_),
	.B1(FE_OFN33_n_1381),
	.Q(n_2009));
   AOI22_X1_50_SVT g79216__1617 (.A0(DPATH_RF_MEMORY_9__6_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__6_),
	.B1(n_1417),
	.Q(n_2008));
   AOI22_X1_50_SVT g79217__2802 (.A0(DPATH_RF_MEMORY_24__4_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__4_),
	.B1(n_1445),
	.Q(n_2007));
   AOI22_X1_50_SVT g79218__1705 (.A0(DPATH_RF_MEMORY_12__6_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__6_),
	.B1(FE_OFN40_n_1391),
	.Q(n_2006));
   AOI22_X1_50_SVT g79219__5122 (.A0(DPATH_RF_MEMORY_28__4_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__4_),
	.B1(FE_OFN31_n_1379),
	.Q(n_2005));
   AOI22_X1_50_SVT g79220__8246 (.A0(DPATH_RF_MEMORY_25__4_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__4_),
	.B1(n_1389),
	.Q(n_2004));
   AOI22_X1_50_SVT g79221__7098 (.A0(DPATH_RF_MEMORY_16__6_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__6_),
	.B1(FE_OFN62_n_1429),
	.Q(n_2003));
   AOI22_X1_50_SVT g79222__6131 (.A0(DPATH_RF_MEMORY_5__4_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__4_),
	.B1(FE_OFN49_n_1404),
	.Q(n_2002));
   AOI22_X1_50_SVT g79223__1881 (.A0(DPATH_RF_MEMORY_1__4_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__4_),
	.B1(n_1434),
	.Q(n_2001));
   AO22_X0_50_SVT g79224__5115 (.A0(DPATH_RF_MEMORY_4__4_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__4_),
	.B1(n_1446),
	.Q(n_2000));
   AOI22_X1_50_SVT g79225__7482 (.A0(DPATH_RF_MEMORY_29__19_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__19_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1999));
   AOI22_X1_50_SVT g79226__4733 (.A0(DPATH_RF_MEMORY_5__26_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__26_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1998));
   AOI22_X1_50_SVT g79227__6161 (.A0(DPATH_RF_MEMORY_1__3_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__3_),
	.B1(n_1434),
	.Q(n_1997));
   AOI22_X1_50_SVT g79228__9315 (.A0(DPATH_RF_MEMORY_8__3_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__3_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1996));
   AOI22_X1_50_SVT g79229__9945 (.A0(DPATH_RF_MEMORY_5__3_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__3_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1995));
   AOI22_X1_50_SVT g79230__2883 (.A0(DPATH_RF_MEMORY_4__3_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__3_),
	.B1(n_1446),
	.Q(n_1994));
   AOI22_X1_50_SVT g79231__2346 (.A0(DPATH_RF_MEMORY_1__6_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__6_),
	.B1(n_1427),
	.Q(n_1993));
   AOI22_X1_50_SVT g79232__1666 (.A0(DPATH_RF_MEMORY_25__3_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__3_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1992));
   AOI22_X1_50_SVT g79233__7410 (.A0(DPATH_RF_MEMORY_28__19_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__19_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1991));
   AOI22_X1_50_SVT g79234__6417 (.A0(DPATH_RF_MEMORY_28__3_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__3_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1990));
   AOI22_X1_50_SVT g79235__5477 (.A0(DPATH_RF_MEMORY_5__6_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__6_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1989));
   AOI22_X1_50_SVT g79236__2398 (.A0(DPATH_RF_MEMORY_24__3_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__3_),
	.B1(n_1445),
	.Q(n_1988));
   AOI22_X1_50_SVT g79237__5107 (.A0(DPATH_RF_MEMORY_8__6_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__6_),
	.B1(n_1403),
	.Q(n_1987));
   AOI22_X1_50_SVT g79238__6260 (.A0(DPATH_RF_MEMORY_20__3_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_19__3_),
	.B1(n_1440),
	.Q(n_1986));
   AOI22_X1_50_SVT g79239__4319 (.A0(DPATH_RF_MEMORY_21__3_),
	.A1(n_1436),
	.B0(DPATH_RF_MEMORY_22__3_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1985));
   AOI22_X1_50_SVT g79240__8428 (.A0(DPATH_RF_MEMORY_9__3_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__3_),
	.B1(n_1399),
	.Q(n_1984));
   AOI22_X1_50_SVT g79241__5526 (.A0(DPATH_RF_MEMORY_12__30_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__30_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1983));
   AOI22_X1_50_SVT g79242__6783 (.A0(DPATH_RF_MEMORY_21__6_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__6_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1982));
   AOI22_X1_50_SVT g79243__3680 (.A0(DPATH_RF_MEMORY_1__26_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__26_),
	.B1(n_1427),
	.Q(n_1981));
   AOI22_X1_50_SVT g79244__1617 (.A0(DPATH_RF_MEMORY_21__29_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__29_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1980));
   AOI22_X1_50_SVT g79245__2802 (.A0(DPATH_RF_MEMORY_12__19_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__19_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1979));
   AOI22_X1_50_SVT g79246__1705 (.A0(DPATH_RF_MEMORY_17__2_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_19__2_),
	.B1(n_1440),
	.Q(n_1978));
   AOI22_X1_50_SVT g79247__5122 (.A0(DPATH_RF_MEMORY_17__6_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_31__6_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1977));
   AOI22_X1_50_SVT g79248__8246 (.A0(DPATH_RF_MEMORY_16__2_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__2_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1976));
   AOI22_X1_50_SVT g79249__7098 (.A0(DPATH_RF_MEMORY_12__2_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__2_),
	.B1(n_1450),
	.Q(n_1975));
   AOI22_X1_50_SVT g79250__6131 (.A0(DPATH_RF_MEMORY_9__2_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__2_),
	.B1(n_1399),
	.Q(n_1974));
   AOI22_X1_50_SVT g79251__1881 (.A0(DPATH_RF_MEMORY_9__19_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__19_),
	.B1(n_1417),
	.Q(n_1973));
   AOI22_X1_50_SVT g79252__5115 (.A0(DPATH_RF_MEMORY_29__2_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__2_),
	.B1(n_1378),
	.Q(n_1972));
   AOI22_X1_50_SVT g79253__7482 (.A0(DPATH_RF_MEMORY_24__2_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__2_),
	.B1(n_1445),
	.Q(n_1971));
   AOI22_X1_50_SVT g79254__4733 (.A0(DPATH_RF_MEMORY_17__25_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_19__25_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1970));
   AOI22_X1_50_SVT g79255__6161 (.A0(DPATH_RF_MEMORY_4__2_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__2_),
	.B1(n_1446),
	.Q(n_1969));
   AOI22_X1_50_SVT g79256__9315 (.A0(DPATH_RF_MEMORY_5__2_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__2_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1968));
   AOI22_X1_50_SVT g79257__9945 (.A0(DPATH_RF_MEMORY_8__2_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__2_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1967));
   AOI22_X1_50_SVT g79258__2883 (.A0(DPATH_RF_MEMORY_29__9_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__9_),
	.B1(n_1378),
	.Q(n_1966));
   AO22_X0_50_SVT g79259__2346 (.A0(DPATH_RF_MEMORY_25__6_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__6_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1965));
   AOI22_X1_50_SVT g79260__1666 (.A0(DPATH_RF_MEMORY_17__1_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_19__1_),
	.B1(n_1440),
	.Q(n_1964));
   AO22_X0_50_SVT g79261__7410 (.A0(DPATH_RF_MEMORY_16__19_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__19_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1963));
   AOI22_X1_50_SVT g79262__6417 (.A0(DPATH_RF_MEMORY_17__5_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_19__5_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1962));
   AOI22_X1_50_SVT g79263__5477 (.A0(DPATH_RF_MEMORY_16__1_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__1_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1961));
   AOI22_X1_50_SVT g79264__2398 (.A0(DPATH_RF_MEMORY_13__1_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__1_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1960));
   AOI22_X1_50_SVT g79265__5107 (.A0(DPATH_RF_MEMORY_12__1_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__1_),
	.B1(n_1450),
	.Q(n_1959));
   AOI22_X1_50_SVT g79266__6260 (.A0(DPATH_RF_MEMORY_29__1_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__1_),
	.B1(n_1378),
	.Q(n_1958));
   AOI22_X1_50_SVT g79267__4319 (.A0(DPATH_RF_MEMORY_24__1_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__1_),
	.B1(n_1445),
	.Q(n_1957));
   AO22_X0_50_SVT g79268__8428 (.A0(DPATH_RF_MEMORY_28__1_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__1_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1956));
   AOI22_X1_50_SVT g79269__5526 (.A0(DPATH_RF_MEMORY_8__19_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__19_),
	.B1(n_1403),
	.Q(n_1955));
   AOI22_X1_50_SVT g79270__6783 (.A0(DPATH_RF_MEMORY_28__5_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__5_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1954));
   AOI22_X1_50_SVT g79271__3680 (.A0(DPATH_RF_MEMORY_5__1_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__1_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1953));
   AOI22_X1_50_SVT g79272__1617 (.A0(DPATH_RF_MEMORY_8__1_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__1_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1952));
   AOI22_X1_50_SVT g79273__2802 (.A0(DPATH_RF_MEMORY_24__5_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__5_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1951));
   AOI22_X1_50_SVT g79274__1705 (.A0(DPATH_RF_MEMORY_5__0_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__0_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1950));
   AOI22_X1_50_SVT g79275__5122 (.A0(DPATH_RF_MEMORY_8__0_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__0_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1949));
   AOI22_X1_50_SVT g79276__8246 (.A0(DPATH_RF_MEMORY_5__19_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__19_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1948));
   AOI22_X1_50_SVT g79277__7098 (.A0(DPATH_RF_MEMORY_4__0_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__0_),
	.B1(n_1446),
	.Q(n_1947));
   AOI22_X1_50_SVT g79278__6131 (.A0(DPATH_RF_MEMORY_29__5_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__5_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1946));
   AOI22_X1_50_SVT g79279__1881 (.A0(DPATH_RF_MEMORY_1__0_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__0_),
	.B1(n_1434),
	.Q(n_1945));
   AOI22_X1_50_SVT g79280__5115 (.A0(DPATH_RF_MEMORY_25__0_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__0_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1944));
   AOI22_X1_50_SVT g79281__7482 (.A0(DPATH_RF_MEMORY_25__5_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__5_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1943));
   AOI22_X1_50_SVT g79282__4733 (.A0(DPATH_RF_MEMORY_29__0_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__0_),
	.B1(n_1378),
	.Q(n_1942));
   AOI22_X1_50_SVT g79283__6161 (.A0(DPATH_RF_MEMORY_28__0_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__0_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1941));
   AOI22_X1_50_SVT g79284__9315 (.A0(DPATH_RF_MEMORY_17__0_),
	.A1(n_1371),
	.B0(DPATH_RF_MEMORY_31__0_),
	.B1(n_1386),
	.Q(n_1940));
   AOI22_X1_50_SVT g79285__9945 (.A0(DPATH_RF_MEMORY_1__19_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__19_),
	.B1(n_1427),
	.Q(n_1939));
   AOI22_X1_50_SVT g79286__2883 (.A0(DPATH_RF_MEMORY_12__5_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__5_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1938));
   AOI22_X1_50_SVT g79287__2346 (.A0(DPATH_RF_MEMORY_20__0_),
	.A1(n_1408),
	.B0(DPATH_RF_MEMORY_19__0_),
	.B1(n_1440),
	.Q(n_1937));
   AOI22_X1_50_SVT g79288__1666 (.A0(DPATH_RF_MEMORY_13__0_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__0_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1936));
   AOI22_X1_50_SVT g79289__7410 (.A0(DPATH_RF_MEMORY_12__0_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__0_),
	.B1(n_1450),
	.Q(n_1935));
   AOI22_X1_50_SVT g79290__6417 (.A0(DPATH_RF_MEMORY_29__29_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__29_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1934));
   AOI22_X1_50_SVT g79291__5477 (.A0(DPATH_RF_MEMORY_9__5_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__5_),
	.B1(n_1417),
	.Q(n_1933));
   AO22_X0_50_SVT g79292__2398 (.A0(DPATH_RF_MEMORY_16__0_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__0_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1932));
   AOI22_X1_50_SVT g79293__5107 (.A0(DPATH_RF_MEMORY_29__25_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__25_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1931));
   AOI22_X1_50_SVT g79294__6260 (.A0(DPATH_RF_MEMORY_16__30_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__30_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1930));
   AOI22_X1_50_SVT g79295__4319 (.A0(DPATH_RF_MEMORY_21__18_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_31__18_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1929));
   AO22_X0_50_SVT g79296__8428 (.A0(DPATH_RF_MEMORY_16__5_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__5_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1928));
   AOI22_X1_50_SVT g79297__5526 (.A0(DPATH_RF_MEMORY_1__5_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__5_),
	.B1(n_1427),
	.Q(n_1927));
   AOI22_X1_50_SVT g79298__6783 (.A0(DPATH_RF_MEMORY_24__25_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__25_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1926));
   AOI22_X1_50_SVT g79299__3680 (.A0(DPATH_RF_MEMORY_4__5_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__5_),
	.B1(n_1420),
	.Q(n_1925));
   AOI22_X1_50_SVT g79300__1617 (.A0(DPATH_RF_MEMORY_25__4_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__4_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1924));
   AOI22_X1_50_SVT g79301__2802 (.A0(DPATH_RF_MEMORY_28__25_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__25_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1923));
   AOI22_X1_50_SVT g79302__1705 (.A0(DPATH_RF_MEMORY_12__18_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__18_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1922));
   AOI22_X1_50_SVT g79303__5122 (.A0(DPATH_RF_MEMORY_13__4_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__4_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1921));
   AO22_X0_50_SVT g79304__8246 (.A0(DPATH_RF_MEMORY_28__29_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__29_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1920));
   AOI22_X1_50_SVT g79305__7098 (.A0(DPATH_RF_MEMORY_9__18_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__18_),
	.B1(n_1417),
	.Q(n_1919));
   AOI22_X1_50_SVT g79306__6131 (.A0(DPATH_RF_MEMORY_24__4_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__4_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1918));
   AOI22_X1_50_SVT g79307__1881 (.A0(DPATH_RF_MEMORY_29__4_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__4_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1917));
   AOI22_X1_50_SVT g79308__5115 (.A0(DPATH_RF_MEMORY_28__4_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__4_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1916));
   AOI22_X1_50_SVT g79309__7482 (.A0(DPATH_RF_MEMORY_16__18_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__18_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1915));
   AOI22_X1_50_SVT g79310__4733 (.A0(DPATH_RF_MEMORY_25__25_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__25_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1914));
   AOI22_X1_50_SVT g79311__6161 (.A0(DPATH_RF_MEMORY_16__4_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__4_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1913));
   AOI22_X1_50_SVT g79312__9315 (.A0(DPATH_RF_MEMORY_29__18_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__18_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1912));
   AOI22_X1_50_SVT g79313__9945 (.A0(DPATH_RF_MEMORY_13__4_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__4_),
	.B1(n_1412),
	.Q(n_1911));
   AOI22_X1_50_SVT g79314__2883 (.A0(DPATH_RF_MEMORY_9__4_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__4_),
	.B1(n_1399),
	.Q(n_1910));
   AOI22_X1_50_SVT g79315__2346 (.A0(DPATH_RF_MEMORY_13__30_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__30_),
	.B1(n_1412),
	.Q(n_1909));
   AOI22_X1_50_SVT g79316__1666 (.A0(DPATH_RF_MEMORY_12__4_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__4_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1908));
   AOI22_X1_50_SVT g79317__7410 (.A0(DPATH_RF_MEMORY_25__18_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__18_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1907));
   AOI22_X1_50_SVT g79318__6417 (.A0(DPATH_RF_MEMORY_16__25_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__25_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1906));
   AOI22_X1_50_SVT g79319__5477 (.A0(DPATH_RF_MEMORY_4__4_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__4_),
	.B1(n_1420),
	.Q(n_1905));
   AO22_X0_50_SVT g79320__2398 (.A0(DPATH_RF_MEMORY_28__18_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__18_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1904));
   AOI22_X1_50_SVT g79321__5107 (.A0(DPATH_RF_MEMORY_8__4_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__4_),
	.B1(n_1403),
	.Q(n_1903));
   AOI22_X1_50_SVT g79322__6260 (.A0(DPATH_RF_MEMORY_1__4_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__4_),
	.B1(n_1427),
	.Q(n_1902));
   AOI22_X1_50_SVT g79323__4319 (.A0(DPATH_RF_MEMORY_16__3_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__3_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1901));
   AOI22_X1_50_SVT g79324__8428 (.A0(DPATH_RF_MEMORY_9__25_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__25_),
	.B1(n_1417),
	.Q(n_1900));
   AOI22_X1_50_SVT g79325__5526 (.A0(DPATH_RF_MEMORY_12__3_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__3_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1899));
   AOI22_X1_50_SVT g79326__6783 (.A0(DPATH_RF_MEMORY_13__3_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__3_),
	.B1(n_1412),
	.Q(n_1898));
   AOI22_X1_50_SVT g79327__3680 (.A0(DPATH_RF_MEMORY_17__28_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__28_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1897));
   AOI22_X1_50_SVT g79328__1617 (.A0(DPATH_RF_MEMORY_1__18_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__18_),
	.B1(n_1427),
	.Q(n_1896));
   AOI22_X1_50_SVT g79329__2802 (.A0(DPATH_RF_MEMORY_9__3_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__3_),
	.B1(n_1417),
	.Q(n_1895));
   AO22_X0_50_SVT g79330__1705 (.A0(DPATH_RF_MEMORY_13__25_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__25_),
	.B1(n_1412),
	.Q(n_1894));
   AOI22_X1_50_SVT g79331__5122 (.A0(DPATH_RF_MEMORY_5__18_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__18_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1893));
   AOI22_X1_50_SVT g79332__8246 (.A0(DPATH_RF_MEMORY_4__3_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__3_),
	.B1(n_1420),
	.Q(n_1892));
   AOI22_X1_50_SVT g79333__7098 (.A0(DPATH_RF_MEMORY_8__3_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__3_),
	.B1(n_1403),
	.Q(n_1891));
   AOI22_X1_50_SVT g79334__6131 (.A0(DPATH_RF_MEMORY_4__18_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__18_),
	.B1(n_1420),
	.Q(n_1890));
   AOI22_X1_50_SVT g79335__1881 (.A0(DPATH_RF_MEMORY_1__3_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__3_),
	.B1(n_1427),
	.Q(n_1889));
   AOI22_X1_50_SVT g79336__5115 (.A0(DPATH_RF_MEMORY_9__30_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__30_),
	.B1(n_1417),
	.Q(n_1888));
   AOI22_X1_50_SVT g79337__7482 (.A0(DPATH_RF_MEMORY_17__3_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_31__3_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1887));
   AOI22_X1_50_SVT g79338__4733 (.A0(DPATH_RF_MEMORY_13__31_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__31_),
	.B1(n_1412),
	.Q(n_1886));
   AOI22_X1_50_SVT g79339__6161 (.A0(DPATH_RF_MEMORY_18__17_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_22__17_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1885));
   AOI22_X1_50_SVT g79340__9315 (.A0(DPATH_RF_MEMORY_21__3_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__3_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1884));
   AOI22_X1_50_SVT g79341__9945 (.A0(DPATH_RF_MEMORY_24__3_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__3_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1883));
   AOI22_X1_50_SVT g79342__2883 (.A0(DPATH_RF_MEMORY_29__3_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__3_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1882));
   AO22_X0_50_SVT g79343__2346 (.A0(DPATH_RF_MEMORY_28__3_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__3_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1881));
   AOI22_X1_50_SVT g79344__1666 (.A0(DPATH_RF_MEMORY_5__25_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__25_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1880));
   AOI22_X1_50_SVT g79345__7410 (.A0(DPATH_RF_MEMORY_20__28_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__28_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1879));
   AOI22_X1_50_SVT g79346__6417 (.A0(DPATH_RF_MEMORY_13__17_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__17_),
	.B1(n_1412),
	.Q(n_1878));
   AOI22_X1_50_SVT g79347__5477 (.A0(DPATH_RF_MEMORY_12__2_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__2_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1877));
   AOI22_X1_50_SVT g79348__2398 (.A0(DPATH_RF_MEMORY_12__17_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__17_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1876));
   AOI22_X1_50_SVT g79349__5107 (.A0(DPATH_RF_MEMORY_9__2_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__2_),
	.B1(n_1417),
	.Q(n_1875));
   AOI22_X1_50_SVT g79350__6260 (.A0(DPATH_RF_MEMORY_13__2_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__2_),
	.B1(n_1412),
	.Q(n_1874));
   AOI22_X1_50_SVT g79351__4319 (.A0(DPATH_RF_MEMORY_16__2_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__2_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1873));
   AOI22_X1_50_SVT g79352__8428 (.A0(DPATH_RF_MEMORY_8__25_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__25_),
	.B1(n_1403),
	.Q(n_1872));
   AOI22_X1_50_SVT g79353__5526 (.A0(DPATH_RF_MEMORY_16__17_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__17_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1871));
   AOI22_X1_50_SVT g79354__6783 (.A0(DPATH_RF_MEMORY_24__6_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__6_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1870));
   AOI22_X1_50_SVT g79355__3680 (.A0(DPATH_RF_MEMORY_9__17_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__17_),
	.B1(n_1417),
	.Q(n_1869));
   AOI22_X1_50_SVT g79356__1617 (.A0(DPATH_RF_MEMORY_4__2_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__2_),
	.B1(n_1420),
	.Q(n_1868));
   AOI22_X1_50_SVT g79357__2802 (.A0(DPATH_RF_MEMORY_8__2_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__2_),
	.B1(n_1403),
	.Q(n_1867));
   AOI22_X1_50_SVT g79358__1705 (.A0(DPATH_RF_MEMORY_1__2_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__2_),
	.B1(n_1427),
	.Q(n_1866));
   AOI22_X1_50_SVT g79359__5122 (.A0(DPATH_RF_MEMORY_21__2_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__2_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1865));
   AOI22_X1_50_SVT g79360__8246 (.A0(DPATH_RF_MEMORY_1__25_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__25_),
	.B1(n_1427),
	.Q(n_1864));
   AOI22_X1_50_SVT g79361__7098 (.A0(DPATH_RF_MEMORY_25__22_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__22_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1863));
   AOI22_X1_50_SVT g79362__6131 (.A0(DPATH_RF_MEMORY_25__17_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__17_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1862));
   AOI22_X1_50_SVT g79363__1881 (.A0(DPATH_RF_MEMORY_18__2_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__2_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1861));
   AOI22_X1_50_SVT g79364__5115 (.A0(DPATH_RF_MEMORY_29__17_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__17_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1860));
   AOI22_X1_50_SVT g79365__7482 (.A0(DPATH_RF_MEMORY_28__2_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__2_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1859));
   AOI22_X1_50_SVT g79366__4733 (.A0(DPATH_RF_MEMORY_25__2_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__2_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1858));
   AO22_X0_50_SVT g79367__6161 (.A0(DPATH_RF_MEMORY_28__17_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__17_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1857));
   AO22_X0_50_SVT g79368__9315 (.A0(DPATH_RF_MEMORY_24__2_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__2_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1856));
   AOI22_X1_50_SVT g79369__9945 (.A0(DPATH_RF_MEMORY_5__24_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__24_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1855));
   AOI22_X1_50_SVT g79370__2883 (.A0(DPATH_RF_MEMORY_17__1_),
	.A1(n_1415),
	.B0(DPATH_RF_MEMORY_18__1_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1854));
   AOI22_X1_50_SVT g79371__2346 (.A0(DPATH_RF_MEMORY_25__28_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__28_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1853));
   AOI22_X1_50_SVT g79372__1666 (.A0(DPATH_RF_MEMORY_20__1_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__1_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1852));
   AOI22_X1_50_SVT g79373__7410 (.A0(DPATH_RF_MEMORY_1__24_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__24_),
	.B1(n_1427),
	.Q(n_1851));
   AOI22_X1_50_SVT g79374__6417 (.A0(DPATH_RF_MEMORY_8__17_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__17_),
	.B1(n_1403),
	.Q(n_1850));
   AOI22_X1_50_SVT g79375__5477 (.A0(DPATH_RF_MEMORY_25__1_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__1_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1849));
   AOI22_X1_50_SVT g79376__2398 (.A0(DPATH_RF_MEMORY_5__17_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__17_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1848));
   AOI22_X1_50_SVT g79377__5107 (.A0(DPATH_RF_MEMORY_28__1_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__1_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1847));
   AOI22_X1_50_SVT g79378__6260 (.A0(DPATH_RF_MEMORY_8__24_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__24_),
	.B1(n_1403),
	.Q(n_1846));
   AOI22_X1_50_SVT g79379__4319 (.A0(DPATH_RF_MEMORY_29__1_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__1_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1845));
   AOI22_X1_50_SVT g79380__8428 (.A0(DPATH_RF_MEMORY_24__1_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__1_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1844));
   AOI22_X1_50_SVT g79381__5526 (.A0(DPATH_RF_MEMORY_1__17_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__17_),
	.B1(n_1427),
	.Q(n_1843));
   AOI22_X1_50_SVT g79382__6783 (.A0(DPATH_RF_MEMORY_17__16_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__16_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1842));
   AOI22_X1_50_SVT g79383__3680 (.A0(DPATH_RF_MEMORY_4__24_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__24_),
	.B1(n_1420),
	.Q(n_1841));
   AOI22_X1_50_SVT g79384__1617 (.A0(DPATH_RF_MEMORY_5__1_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__1_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1840));
   AOI22_X1_50_SVT g79385__2802 (.A0(DPATH_RF_MEMORY_4__1_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__1_),
	.B1(n_1420),
	.Q(n_1839));
   AOI22_X1_50_SVT g79386__1705 (.A0(DPATH_RF_MEMORY_12__1_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__1_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1838));
   AOI22_X1_50_SVT g79387__5122 (.A0(DPATH_RF_MEMORY_29__28_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__28_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1837));
   AOI22_X1_50_SVT g79388__8246 (.A0(DPATH_RF_MEMORY_12__29_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__29_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1836));
   NAND2_X1_50_SVT g79389__7098 (.A(n_3),
	.B(n_1468),
	.Q(n_2202));
   AOI22_X1_50_SVT g79390__6131 (.A0(DPATH_RF_MEMORY_16__1_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__1_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1835));
   AOI22_X1_50_SVT g79391__1881 (.A0(DPATH_RF_MEMORY_13__1_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__1_),
	.B1(n_1412),
	.Q(n_1834));
   AOI22_X1_50_SVT g79392__5115 (.A0(DPATH_RF_MEMORY_8__30_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__30_),
	.B1(n_1403),
	.Q(n_1833));
   AOI22_X1_50_SVT g79393__7482 (.A0(DPATH_RF_MEMORY_9__1_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__1_),
	.B1(n_1417),
	.Q(n_1832));
   AOI22_X1_50_SVT g79394__4733 (.A0(DPATH_RF_MEMORY_12__0_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__0_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1831));
   AOI22_X1_50_SVT g79395__6161 (.A0(DPATH_RF_MEMORY_9__0_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__0_),
	.B1(n_1417),
	.Q(n_1830));
   AOI22_X1_50_SVT g79396__9315 (.A0(DPATH_RF_MEMORY_25__16_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__16_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1829));
   AO22_X0_50_SVT g79397__9945 (.A0(DPATH_RF_MEMORY_16__0_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__0_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1828));
   AOI22_X1_50_SVT g79398__2883 (.A0(DPATH_RF_MEMORY_28__28_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__28_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1827));
   AOI22_X1_50_SVT g79399__2346 (.A0(DPATH_RF_MEMORY_24__24_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__24_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1826));
   AOI22_X1_50_SVT g79400__1666 (.A0(DPATH_RF_MEMORY_24__16_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__16_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1825));
   AOI22_X1_50_SVT g79401__7410 (.A0(DPATH_RF_MEMORY_20__0_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__0_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1824));
   AOI22_X1_50_SVT g79402__6417 (.A0(DPATH_RF_MEMORY_29__16_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__16_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1823));
   AOI22_X1_50_SVT g79403__5477 (.A0(DPATH_RF_MEMORY_29__24_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__24_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1822));
   AOI22_X1_50_SVT g79404__2398 (.A0(DPATH_RF_MEMORY_5__0_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__0_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1821));
   AOI22_X1_50_SVT g79405__5107 (.A0(DPATH_RF_MEMORY_28__16_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__16_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1820));
   AOI22_X1_50_SVT g79406__6260 (.A0(DPATH_RF_MEMORY_8__0_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__0_),
	.B1(n_1403),
	.Q(n_1819));
   AOI22_X1_50_SVT g79407__4319 (.A0(DPATH_RF_MEMORY_4__0_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__0_),
	.B1(n_1420),
	.Q(n_1818));
   AOI22_X1_50_SVT g79408__8428 (.A0(DPATH_RF_MEMORY_29__31_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__31_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1817));
   AOI22_X1_50_SVT g79409__5526 (.A0(DPATH_RF_MEMORY_28__24_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__24_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1816));
   AOI22_X1_50_SVT g79410__6783 (.A0(DPATH_RF_MEMORY_18__0_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__0_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1815));
   AOI22_X1_50_SVT g79411__3680 (.A0(DPATH_RF_MEMORY_25__0_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__0_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1814));
   AOI22_X1_50_SVT g79412__1617 (.A0(DPATH_RF_MEMORY_24__28_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__28_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1813));
   AOI22_X1_50_SVT g79413__2802 (.A0(DPATH_RF_MEMORY_24__0_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__0_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1812));
   AOI22_X1_50_SVT g79414__1705 (.A0(DPATH_RF_MEMORY_4__16_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__16_),
	.B1(n_1420),
	.Q(n_1811));
   AOI22_X1_50_SVT g79415__5122 (.A0(DPATH_RF_MEMORY_29__0_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__0_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1810));
   AOI22_X1_50_SVT g79416__8246 (.A0(DPATH_RF_MEMORY_1__16_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__16_),
	.B1(n_1427),
	.Q(n_1809));
   AOI22_X1_50_SVT g79417__7098 (.A0(DPATH_RF_MEMORY_28__0_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__0_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1808));
   AOI22_X1_50_SVT g79418__6131 (.A0(DPATH_RF_MEMORY_20__24_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__24_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1807));
   AOI22_X1_50_SVT g79419__1881 (.A0(DPATH_RF_MEMORY_17__31_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_18__31_),
	.B1(FE_OFN63_n_1432),
	.Q(n_1806));
   AOI22_X1_50_SVT g79420__5115 (.A0(DPATH_RF_MEMORY_5__30_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__30_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1805));
   AOI22_X1_50_SVT g79421__7482 (.A0(DPATH_RF_MEMORY_9__16_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__16_),
	.B1(n_1417),
	.Q(n_1804));
   AOI22_X1_50_SVT g79422__4733 (.A0(DPATH_RF_MEMORY_16__16_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__16_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1803));
   AOI22_X1_50_SVT g79423__6161 (.A0(DPATH_RF_MEMORY_20__31_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__31_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1802));
   AOI22_X1_50_SVT g79424__9315 (.A0(DPATH_RF_MEMORY_1__30_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__30_),
	.B1(n_1427),
	.Q(n_1801));
   AOI22_X1_50_SVT g79425__9945 (.A0(DPATH_RF_MEMORY_13__16_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__16_),
	.B1(n_1412),
	.Q(n_1800));
   AOI22_X1_50_SVT g79426__2883 (.A0(DPATH_RF_MEMORY_29__31_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__31_),
	.B1(n_1378),
	.Q(n_1799));
   AOI22_X1_50_SVT g79427__2346 (.A0(DPATH_RF_MEMORY_12__16_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__16_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1798));
   AOI22_X1_50_SVT g79428__1666 (.A0(DPATH_RF_MEMORY_24__31_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__31_),
	.B1(n_1445),
	.Q(n_1797));
   AOI22_X1_50_SVT g79429__7410 (.A0(DPATH_RF_MEMORY_21__24_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__24_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1796));
   AOI22_X1_50_SVT g79430__6417 (.A0(DPATH_RF_MEMORY_13__15_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__15_),
	.B1(n_1412),
	.Q(n_1795));
   AOI22_X1_50_SVT g79431__5477 (.A0(DPATH_RF_MEMORY_28__31_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__31_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1794));
   AOI22_X1_50_SVT g79432__2398 (.A0(DPATH_RF_MEMORY_25__31_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__31_),
	.B1(n_1389),
	.Q(n_1793));
   AOI22_X1_50_SVT g79433__5107 (.A0(DPATH_RF_MEMORY_12__24_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__24_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1792));
   AOI22_X1_50_SVT g79434__6260 (.A0(DPATH_RF_MEMORY_16__15_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__15_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1791));
   AOI22_X1_50_SVT g79435__4319 (.A0(DPATH_RF_MEMORY_5__31_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__31_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1790));
   AOI22_X1_50_SVT g79436__8428 (.A0(DPATH_RF_MEMORY_4__31_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__31_),
	.B1(n_1446),
	.Q(n_1789));
   AO22_X0_50_SVT g79437__5526 (.A0(DPATH_RF_MEMORY_9__15_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__15_),
	.B1(n_1417),
	.Q(n_1788));
   AOI22_X1_50_SVT g79438__6783 (.A0(DPATH_RF_MEMORY_13__31_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__31_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1787));
   AOI22_X1_50_SVT g79439__3680 (.A0(DPATH_RF_MEMORY_8__24_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__24_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1786));
   AOI22_X1_50_SVT g79440__1617 (.A0(DPATH_RF_MEMORY_9__24_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__24_),
	.B1(n_1417),
	.Q(n_1785));
   AOI22_X1_50_SVT g79441__2802 (.A0(DPATH_RF_MEMORY_16__31_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__31_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1784));
   AOI22_X1_50_SVT g79442__1705 (.A0(DPATH_RF_MEMORY_12__31_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__31_),
	.B1(n_1450),
	.Q(n_1783));
   AOI22_X1_50_SVT g79443__5122 (.A0(DPATH_RF_MEMORY_9__31_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__31_),
	.B1(n_1399),
	.Q(n_1782));
   AOI22_X1_50_SVT g79444__8246 (.A0(DPATH_RF_MEMORY_5__28_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__28_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1781));
   AOI22_X1_50_SVT g79445__7098 (.A0(DPATH_RF_MEMORY_21__15_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__15_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1780));
   AOI22_X1_50_SVT g79446__6131 (.A0(DPATH_RF_MEMORY_16__30_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__30_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1779));
   AOI22_X1_50_SVT g79447__1881 (.A0(DPATH_RF_MEMORY_9__30_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__30_),
	.B1(n_1399),
	.Q(n_1778));
   AOI22_X1_50_SVT g79448__5115 (.A0(DPATH_RF_MEMORY_13__30_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__30_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1777));
   AOI22_X1_50_SVT g79449__7482 (.A0(DPATH_RF_MEMORY_12__30_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__30_),
	.B1(n_1450),
	.Q(n_1776));
   AOI22_X1_50_SVT g79450__4733 (.A0(DPATH_RF_MEMORY_1__30_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__30_),
	.B1(n_1434),
	.Q(n_1775));
   AOI22_X1_50_SVT g79451__6161 (.A0(DPATH_RF_MEMORY_8__28_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__28_),
	.B1(n_1403),
	.Q(n_1774));
   AO22_X0_50_SVT g79452 (.A0(DPATH_RF_MEMORY_16__24_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__24_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1773));
   AOI22_X1_50_SVT g79453 (.A0(DPATH_RF_MEMORY_8__15_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__15_),
	.B1(n_1403),
	.Q(n_1772));
   AOI22_X1_50_SVT g79454 (.A0(DPATH_RF_MEMORY_8__30_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__30_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1771));
   AOI22_X1_50_SVT g79455 (.A0(DPATH_RF_MEMORY_4__30_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__30_),
	.B1(n_1446),
	.Q(n_1770));
   AOI22_X1_50_SVT g79456 (.A0(DPATH_RF_MEMORY_20__30_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__30_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1769));
   AOI22_X1_50_SVT g79457 (.A0(DPATH_RF_MEMORY_4__15_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__15_),
	.B1(n_1420),
	.Q(n_1768));
   AOI22_X1_50_SVT g79458 (.A0(DPATH_RF_MEMORY_21__30_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__30_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1767));
   AOI22_X1_50_SVT g79459 (.A0(DPATH_RF_MEMORY_24__30_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__30_),
	.B1(n_1445),
	.Q(n_1766));
   AOI22_X1_50_SVT g79460 (.A0(DPATH_RF_MEMORY_21__30_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__30_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1765));
   AOI22_X1_50_SVT g79461 (.A0(DPATH_RF_MEMORY_1__15_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__15_),
	.B1(n_1427),
	.Q(n_1764));
   AOI22_X1_50_SVT g79462 (.A0(DPATH_RF_MEMORY_25__30_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__30_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1763));
   AO22_X0_50_SVT g79463 (.A0(DPATH_RF_MEMORY_28__30_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__30_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1762));
   AOI22_X1_50_SVT g79464 (.A0(DPATH_RF_MEMORY_18__15_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__15_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1761));
   AOI22_X1_50_SVT g79465 (.A0(DPATH_RF_MEMORY_8__29_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__29_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1760));
   AOI22_X1_50_SVT g79466 (.A0(DPATH_RF_MEMORY_1__29_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__29_),
	.B1(n_1434),
	.Q(n_1759));
   AOI22_X1_50_SVT g79467 (.A0(DPATH_RF_MEMORY_5__29_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__29_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1758));
   AOI22_X1_50_SVT g79468 (.A0(DPATH_RF_MEMORY_4__29_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__29_),
	.B1(n_1446),
	.Q(n_1757));
   AOI22_X1_50_SVT g79469 (.A0(DPATH_RF_MEMORY_28__15_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__15_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1756));
   AOI22_X1_50_SVT g79470 (.A0(DPATH_RF_MEMORY_9__28_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__28_),
	.B1(n_1417),
	.Q(n_1755));
   AOI22_X1_50_SVT g79471 (.A0(DPATH_RF_MEMORY_24__29_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__29_),
	.B1(n_1445),
	.Q(n_1754));
   AOI22_X1_50_SVT g79472 (.A0(DPATH_RF_MEMORY_28__29_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__29_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1753));
   AOI22_X1_50_SVT g79473 (.A0(DPATH_RF_MEMORY_25__29_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__29_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1752));
   AOI22_X1_50_SVT g79474 (.A0(DPATH_RF_MEMORY_29__15_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__15_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1751));
   AOI22_X1_50_SVT g79475 (.A0(DPATH_RF_MEMORY_21__29_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__29_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1750));
   AOI22_X1_50_SVT g79476 (.A0(DPATH_RF_MEMORY_25__15_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__15_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1749));
   AOI22_X1_50_SVT g79477 (.A0(DPATH_RF_MEMORY_20__29_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__29_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1748));
   AOI22_X1_50_SVT g79478 (.A0(DPATH_RF_MEMORY_16__29_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__29_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1747));
   AOI22_X1_50_SVT g79479 (.A0(DPATH_RF_MEMORY_13__23_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__23_),
	.B1(n_1412),
	.Q(n_1746));
   AOI22_X1_50_SVT g79480 (.A0(DPATH_RF_MEMORY_9__29_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__29_),
	.B1(n_1399),
	.Q(n_1745));
   AOI22_X1_50_SVT g79481 (.A0(DPATH_RF_MEMORY_12__23_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__23_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1744));
   AOI22_X1_50_SVT g79482 (.A0(DPATH_RF_MEMORY_24__15_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__15_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1743));
   AO22_X0_50_SVT g79483 (.A0(DPATH_RF_MEMORY_13__29_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__29_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1742));
   AOI22_X1_50_SVT g79484 (.A0(DPATH_RF_MEMORY_12__31_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__31_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1741));
   AOI22_X1_50_SVT g79485 (.A0(DPATH_RF_MEMORY_17__14_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__14_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1740));
   AOI22_X1_50_SVT g79486 (.A0(DPATH_RF_MEMORY_28__28_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__28_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1739));
   AOI22_X1_50_SVT g79487 (.A0(DPATH_RF_MEMORY_25__31_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__31_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1738));
   AOI22_X1_50_SVT g79488 (.A0(DPATH_RF_MEMORY_25__28_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__28_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1737));
   AOI22_X1_50_SVT g79489 (.A0(DPATH_RF_MEMORY_16__28_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__28_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1736));
   AOI22_X1_50_SVT g79490 (.A0(DPATH_RF_MEMORY_16__23_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__23_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1735));
   AOI22_X1_50_SVT g79491 (.A0(DPATH_RF_MEMORY_29__28_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__28_),
	.B1(n_1378),
	.Q(n_1734));
   AOI22_X1_50_SVT g79492 (.A0(DPATH_RF_MEMORY_24__28_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__28_),
	.B1(n_1445),
	.Q(n_1733));
   AOI22_X1_50_SVT g79493 (.A0(DPATH_RF_MEMORY_20__14_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__14_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1732));
   AOI22_X1_50_SVT g79494 (.A0(DPATH_RF_MEMORY_9__23_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__23_),
	.B1(n_1417),
	.Q(n_1731));
   AOI22_X1_50_SVT g79495 (.A0(DPATH_RF_MEMORY_12__28_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__28_),
	.B1(n_1450),
	.Q(n_1730));
   AOI22_X1_50_SVT g79496 (.A0(DPATH_RF_MEMORY_16__28_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__28_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1729));
   AOI22_X1_50_SVT g79497 (.A0(DPATH_RF_MEMORY_9__28_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__28_),
	.B1(n_1399),
	.Q(n_1728));
   AOI22_X1_50_SVT g79498 (.A0(DPATH_RF_MEMORY_13__28_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__28_),
	.B1(n_1412),
	.Q(n_1727));
   AOI22_X1_50_SVT g79499 (.A0(DPATH_RF_MEMORY_4__28_),
	.A1(n_1380),
	.B0(DPATH_RF_MEMORY_3__28_),
	.B1(n_1446),
	.Q(n_1726));
   AOI22_X1_50_SVT g79500 (.A0(DPATH_RF_MEMORY_24__14_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__14_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1725));
   AOI22_X1_50_SVT g79501 (.A0(DPATH_RF_MEMORY_1__28_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__28_),
	.B1(n_1434),
	.Q(n_1724));
   AOI22_X1_50_SVT g79502 (.A0(DPATH_RF_MEMORY_8__28_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__28_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1723));
   AOI22_X1_50_SVT g79503 (.A0(DPATH_RF_MEMORY_28__14_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__14_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1722));
   AOI22_X1_50_SVT g79504 (.A0(DPATH_RF_MEMORY_13__27_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__27_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1721));
   AOI22_X1_50_SVT g79505 (.A0(DPATH_RF_MEMORY_12__27_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__27_),
	.B1(n_1450),
	.Q(n_1720));
   AOI22_X1_50_SVT g79506 (.A0(DPATH_RF_MEMORY_29__14_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__14_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1719));
   AOI22_X1_50_SVT g79507 (.A0(DPATH_RF_MEMORY_16__27_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__27_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1718));
   AOI22_X1_50_SVT g79508 (.A0(DPATH_RF_MEMORY_9__27_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__27_),
	.B1(n_1399),
	.Q(n_1717));
   AOI22_X1_50_SVT g79509 (.A0(DPATH_RF_MEMORY_25__14_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__14_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1716));
   AOI22_X1_50_SVT g79510 (.A0(DPATH_RF_MEMORY_29__27_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__27_),
	.B1(n_1378),
	.Q(n_1715));
   AOI22_X1_50_SVT g79511 (.A0(DPATH_RF_MEMORY_25__27_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__27_),
	.B1(n_1389),
	.Q(n_1714));
   AOI22_X1_50_SVT g79512 (.A0(DPATH_RF_MEMORY_24__27_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__27_),
	.B1(n_1445),
	.Q(n_1713));
   AOI22_X1_50_SVT g79513 (.A0(DPATH_RF_MEMORY_12__28_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__28_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1712));
   AOI22_X1_50_SVT g79514 (.A0(DPATH_RF_MEMORY_29__25_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__25_),
	.B1(n_1378),
	.Q(n_1711));
   AOI22_X1_50_SVT g79515 (.A0(DPATH_RF_MEMORY_4__27_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__27_),
	.B1(n_1446),
	.Q(n_1710));
   AOI22_X1_50_SVT g79516 (.A0(DPATH_RF_MEMORY_8__27_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__27_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1709));
   AOI22_X1_50_SVT g79517 (.A0(DPATH_RF_MEMORY_4__14_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__14_),
	.B1(n_1420),
	.Q(n_1708));
   AOI22_X1_50_SVT g79518 (.A0(DPATH_RF_MEMORY_1__27_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__27_),
	.B1(n_1434),
	.Q(n_1707));
   AOI22_X1_50_SVT g79519 (.A0(DPATH_RF_MEMORY_1__26_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__26_),
	.B1(n_1434),
	.Q(n_1706));
   AOI22_X1_50_SVT g79520 (.A0(DPATH_RF_MEMORY_1__14_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__14_),
	.B1(n_1427),
	.Q(n_1705));
   AOI22_X1_50_SVT g79521 (.A0(DPATH_RF_MEMORY_5__26_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__26_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1704));
   AOI22_X1_50_SVT g79522 (.A0(DPATH_RF_MEMORY_8__26_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__26_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1703));
   AOI22_X1_50_SVT g79523 (.A0(DPATH_RF_MEMORY_4__26_),
	.A1(n_1380),
	.B0(DPATH_RF_MEMORY_3__26_),
	.B1(n_1446),
	.Q(n_1702));
   AOI22_X1_50_SVT g79524 (.A0(DPATH_RF_MEMORY_29__23_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__23_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1701));
   AOI22_X1_50_SVT g79525 (.A0(DPATH_RF_MEMORY_18__30_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__30_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1700));
   AOI22_X1_50_SVT g79526 (.A0(DPATH_RF_MEMORY_16__14_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__14_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1699));
   AOI22_X1_50_SVT g79527 (.A0(DPATH_RF_MEMORY_24__26_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__26_),
	.B1(n_1445),
	.Q(n_1698));
   AOI22_X1_50_SVT g79528 (.A0(DPATH_RF_MEMORY_28__26_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__26_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1697));
   AOI22_X1_50_SVT g79529 (.A0(DPATH_RF_MEMORY_17__27_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__27_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1696));
   AOI22_X1_50_SVT g79530 (.A0(DPATH_RF_MEMORY_12__14_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__14_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1695));
   AOI22_X1_50_SVT g79531 (.A0(DPATH_RF_MEMORY_25__26_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__26_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1694));
   AOI22_X1_50_SVT g79532 (.A0(DPATH_RF_MEMORY_21__26_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__26_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1693));
   AOI22_X1_50_SVT g79533 (.A0(DPATH_RF_MEMORY_25__23_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__23_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1692));
   AOI22_X1_50_SVT g79534 (.A0(DPATH_RF_MEMORY_24__31_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__31_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1691));
   AOI22_X1_50_SVT g79535 (.A0(DPATH_RF_MEMORY_13__14_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__14_),
	.B1(n_1412),
	.Q(n_1690));
   AOI22_X1_50_SVT g79536 (.A0(DPATH_RF_MEMORY_20__26_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__26_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1689));
   AOI22_X1_50_SVT g79537 (.A0(DPATH_RF_MEMORY_13__26_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__26_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1688));
   AOI22_X1_50_SVT g79538 (.A0(DPATH_RF_MEMORY_12__26_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__26_),
	.B1(n_1450),
	.Q(n_1687));
   AOI22_X1_50_SVT g79539 (.A0(DPATH_RF_MEMORY_9__14_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__14_),
	.B1(n_1417),
	.Q(n_1686));
   AO22_X0_50_SVT g79540 (.A0(DPATH_RF_MEMORY_16__26_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__26_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1685));
   AOI22_X1_50_SVT g79541 (.A0(DPATH_RF_MEMORY_17__25_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_19__25_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1684));
   AOI22_X1_50_SVT g79542 (.A0(DPATH_RF_MEMORY_24__23_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__23_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1683));
   AOI22_X1_50_SVT g79543 (.A0(DPATH_RF_MEMORY_4__13_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__13_),
	.B1(n_1420),
	.Q(n_1682));
   AOI22_X1_50_SVT g79544 (.A0(DPATH_RF_MEMORY_25__25_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__25_),
	.B1(n_1389),
	.Q(n_1681));
   AOI22_X1_50_SVT g79545 (.A0(DPATH_RF_MEMORY_24__25_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__25_),
	.B1(n_1445),
	.Q(n_1680));
   AOI22_X1_50_SVT g79546 (.A0(DPATH_RF_MEMORY_28__30_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__30_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1679));
   AOI22_X1_50_SVT g79547 (.A0(DPATH_RF_MEMORY_28__25_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__25_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1678));
   AOI22_X1_50_SVT g79548 (.A0(DPATH_RF_MEMORY_8__13_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__13_),
	.B1(n_1403),
	.Q(n_1677));
   AOI22_X1_50_SVT g79549 (.A0(DPATH_RF_MEMORY_16__25_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__25_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1676));
   AOI22_X1_50_SVT g79550 (.A0(DPATH_RF_MEMORY_5__13_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__13_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1675));
   AOI22_X1_50_SVT g79551 (.A0(DPATH_RF_MEMORY_4__23_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__23_),
	.B1(n_1420),
	.Q(n_1674));
   AOI22_X1_50_SVT g79552 (.A0(DPATH_RF_MEMORY_13__25_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__25_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1673));
   AOI22_X1_50_SVT g79553 (.A0(DPATH_RF_MEMORY_9__25_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__25_),
	.B1(n_1399),
	.Q(n_1672));
   AOI22_X1_50_SVT g79554 (.A0(DPATH_RF_MEMORY_1__13_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__13_),
	.B1(n_1427),
	.Q(n_1671));
   AOI22_X1_50_SVT g79555 (.A0(DPATH_RF_MEMORY_4__25_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__25_),
	.B1(n_1446),
	.Q(n_1670));
   AOI22_X1_50_SVT g79556 (.A0(DPATH_RF_MEMORY_8__25_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__25_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1669));
   AO22_X0_50_SVT g79557 (.A0(DPATH_RF_MEMORY_1__25_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__25_),
	.B1(n_1434),
	.Q(n_1668));
   AOI22_X1_50_SVT g79558 (.A0(DPATH_RF_MEMORY_22__24_),
	.A1(FE_OFN65_n_1438),
	.B0(DPATH_RF_MEMORY_31__24_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1667));
   AOI22_X1_50_SVT g79559 (.A0(DPATH_RF_MEMORY_8__23_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__23_),
	.B1(n_1403),
	.Q(n_1666));
   AOI22_X1_50_SVT g79560 (.A0(DPATH_RF_MEMORY_20__27_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__27_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1665));
   AOI22_X1_50_SVT g79561 (.A0(DPATH_RF_MEMORY_24__24_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__24_),
	.B1(n_1445),
	.Q(n_1664));
   AOI22_X1_50_SVT g79562 (.A0(DPATH_RF_MEMORY_25__24_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__24_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1663));
   AOI22_X1_50_SVT g79563 (.A0(DPATH_RF_MEMORY_29__13_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__13_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1662));
   AOI22_X1_50_SVT g79564 (.A0(DPATH_RF_MEMORY_29__24_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__24_),
	.B1(n_1378),
	.Q(n_1661));
   AOI22_X1_50_SVT g79565 (.A0(DPATH_RF_MEMORY_28__13_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__13_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1660));
   AOI22_X1_50_SVT g79566 (.A0(DPATH_RF_MEMORY_28__24_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__24_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1659));
   AOI22_X1_50_SVT g79567 (.A0(DPATH_RF_MEMORY_1__23_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__23_),
	.B1(n_1427),
	.Q(n_1658));
   AOI22_X1_50_SVT g79568 (.A0(DPATH_RF_MEMORY_25__13_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__13_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1657));
   AOI22_X1_50_SVT g79569 (.A0(DPATH_RF_MEMORY_9__24_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__24_),
	.B1(n_1399),
	.Q(n_1656));
   AOI22_X1_50_SVT g79570 (.A0(DPATH_RF_MEMORY_13__24_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__24_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1655));
   AO22_X0_50_SVT g79571 (.A0(DPATH_RF_MEMORY_16__24_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__24_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1654));
   AOI22_X1_50_SVT g79572 (.A0(DPATH_RF_MEMORY_21__13_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__13_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1653));
   AOI22_X1_50_SVT g79573 (.A0(DPATH_RF_MEMORY_4__24_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__24_),
	.B1(n_1446),
	.Q(n_1652));
   AOI22_X1_50_SVT g79574 (.A0(DPATH_RF_MEMORY_29__30_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__30_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1651));
   AOI22_X1_50_SVT g79575 (.A0(DPATH_RF_MEMORY_5__24_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__24_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1650));
   AOI22_X1_50_SVT g79576 (.A0(DPATH_RF_MEMORY_12__23_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__23_),
	.B1(n_1450),
	.Q(n_1649));
   AOI22_X1_50_SVT g79577 (.A0(DPATH_RF_MEMORY_13__22_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__22_),
	.B1(n_1412),
	.Q(n_1648));
   AOI22_X1_50_SVT g79578 (.A0(DPATH_RF_MEMORY_18__13_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__13_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1647));
   AOI22_X1_50_SVT g79579 (.A0(DPATH_RF_MEMORY_16__23_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__23_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1646));
   AOI22_X1_50_SVT g79580 (.A0(DPATH_RF_MEMORY_13__23_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__23_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1645));
   AOI22_X1_50_SVT g79581 (.A0(DPATH_RF_MEMORY_9__23_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__23_),
	.B1(n_1399),
	.Q(n_1644));
   AOI22_X1_50_SVT g79582 (.A0(DPATH_RF_MEMORY_13__13_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__13_),
	.B1(n_1412),
	.Q(n_1643));
   AOI22_X1_50_SVT g79583 (.A0(DPATH_RF_MEMORY_4__23_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__23_),
	.B1(n_1446),
	.Q(n_1642));
   AOI22_X1_50_SVT g79584 (.A0(DPATH_RF_MEMORY_5__23_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__23_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1641));
   AOI22_X1_50_SVT g79585 (.A0(DPATH_RF_MEMORY_12__22_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__22_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1640));
   AOI22_X1_50_SVT g79586 (.A0(DPATH_RF_MEMORY_1__23_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__23_),
	.B1(n_1434),
	.Q(n_1639));
   AOI22_X1_50_SVT g79587 (.A0(DPATH_RF_MEMORY_16__13_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__13_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1638));
   AOI22_X1_50_SVT g79588 (.A0(DPATH_RF_MEMORY_29__27_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__27_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1637));
   AOI22_X1_50_SVT g79589 (.A0(DPATH_RF_MEMORY_20__23_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__23_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1636));
   AOI22_X1_50_SVT g79590 (.A0(DPATH_RF_MEMORY_21__23_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__23_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1635));
   AOI22_X1_50_SVT g79591 (.A0(DPATH_RF_MEMORY_25__23_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__23_),
	.B1(n_1389),
	.Q(n_1634));
   AOI22_X1_50_SVT g79592 (.A0(DPATH_RF_MEMORY_16__22_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__22_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1633));
   AOI22_X1_50_SVT g79593 (.A0(DPATH_RF_MEMORY_29__23_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__23_),
	.B1(n_1378),
	.Q(n_1632));
   AO22_X0_50_SVT g79594 (.A0(DPATH_RF_MEMORY_9__13_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__13_),
	.B1(n_1417),
	.Q(n_1631));
   AOI22_X1_50_SVT g79595 (.A0(DPATH_RF_MEMORY_8__5_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__5_),
	.B1(n_1403),
	.Q(n_1630));
   AO22_X0_50_SVT g79596 (.A0(DPATH_RF_MEMORY_24__23_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__23_),
	.B1(n_1445),
	.Q(n_1629));
   AOI22_X1_50_SVT g79597 (.A0(DPATH_RF_MEMORY_9__22_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__22_),
	.B1(n_1417),
	.Q(n_1628));
   AOI22_X1_50_SVT g79598 (.A0(DPATH_RF_MEMORY_4__22_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__22_),
	.B1(n_1446),
	.Q(n_1627));
   AOI22_X1_50_SVT g79599 (.A0(DPATH_RF_MEMORY_16__12_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__12_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1626));
   AOI22_X1_50_SVT g79600 (.A0(DPATH_RF_MEMORY_8__22_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__22_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1625));
   AOI22_X1_50_SVT g79601 (.A0(DPATH_RF_MEMORY_9__31_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__31_),
	.B1(n_1417),
	.Q(n_1624));
   AOI22_X1_50_SVT g79602 (.A0(DPATH_RF_MEMORY_5__22_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__22_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1623));
   AOI22_X1_50_SVT g79603 (.A0(DPATH_RF_MEMORY_1__22_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__22_),
	.B1(n_1434),
	.Q(n_1622));
   AOI22_X1_50_SVT g79604 (.A0(DPATH_RF_MEMORY_9__12_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__12_),
	.B1(n_1417),
	.Q(n_1621));
   AOI22_X1_50_SVT g79605 (.A0(DPATH_RF_MEMORY_24__22_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__22_),
	.B1(n_1445),
	.Q(n_1620));
   AOI22_X1_50_SVT g79606 (.A0(DPATH_RF_MEMORY_28__27_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__27_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1619));
   AOI22_X1_50_SVT g79607 (.A0(DPATH_RF_MEMORY_29__22_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__22_),
	.B1(n_1378),
	.Q(n_1618));
   AO22_X0_50_SVT g79608 (.A0(DPATH_RF_MEMORY_25__30_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__30_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1617));
   AO22_X0_50_SVT g79609 (.A0(DPATH_RF_MEMORY_13__12_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__12_),
	.B1(n_1412),
	.Q(n_1616));
   AOI22_X1_50_SVT g79610 (.A0(DPATH_RF_MEMORY_16__31_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__31_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1615));
   AOI22_X1_50_SVT g79611 (.A0(DPATH_RF_MEMORY_17__22_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__22_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1614));
   AOI22_X1_50_SVT g79612 (.A0(DPATH_RF_MEMORY_20__22_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__22_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1613));
   AOI22_X1_50_SVT g79613 (.A0(DPATH_RF_MEMORY_12__22_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__22_),
	.B1(n_1450),
	.Q(n_1612));
   AOI22_X1_50_SVT g79614 (.A0(DPATH_RF_MEMORY_9__22_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__22_),
	.B1(n_1399),
	.Q(n_1611));
   AO22_X0_50_SVT g79615 (.A0(DPATH_RF_MEMORY_16__22_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__22_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1610));
   AOI22_X1_50_SVT g79616 (.A0(DPATH_RF_MEMORY_4__22_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__22_),
	.B1(n_1420),
	.Q(n_1609));
   AOI22_X1_50_SVT g79617 (.A0(DPATH_RF_MEMORY_8__21_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__21_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1608));
   AOI22_X1_50_SVT g79618 (.A0(DPATH_RF_MEMORY_21__12_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__12_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1607));
   AOI22_X1_50_SVT g79619 (.A0(DPATH_RF_MEMORY_1__21_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__21_),
	.B1(n_1434),
	.Q(n_1606));
   AOI22_X1_50_SVT g79620 (.A0(DPATH_RF_MEMORY_5__21_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__21_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1605));
   AOI22_X1_50_SVT g79621 (.A0(DPATH_RF_MEMORY_4__21_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__21_),
	.B1(n_1446),
	.Q(n_1604));
   AOI22_X1_50_SVT g79622 (.A0(DPATH_RF_MEMORY_25__27_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__27_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1603));
   AOI22_X1_50_SVT g79623 (.A0(DPATH_RF_MEMORY_24__21_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__21_),
	.B1(n_1445),
	.Q(n_1602));
   AOI22_X1_50_SVT g79624 (.A0(DPATH_RF_MEMORY_8__12_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__12_),
	.B1(n_1403),
	.Q(n_1601));
   AOI22_X1_50_SVT g79625 (.A0(DPATH_RF_MEMORY_28__21_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__21_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1600));
   AOI22_X1_50_SVT g79626 (.A0(DPATH_RF_MEMORY_25__21_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__21_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1599));
   AOI22_X1_50_SVT g79627 (.A0(DPATH_RF_MEMORY_8__22_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__22_),
	.B1(n_1403),
	.Q(n_1598));
   AOI22_X1_50_SVT g79628 (.A0(DPATH_RF_MEMORY_17__21_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__21_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1597));
   AOI22_X1_50_SVT g79629 (.A0(DPATH_RF_MEMORY_1__22_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__22_),
	.B1(n_1427),
	.Q(n_1596));
   AOI22_X1_50_SVT g79630 (.A0(DPATH_RF_MEMORY_5__12_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__12_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1595));
   AOI22_X1_50_SVT g79631 (.A0(DPATH_RF_MEMORY_21__21_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__21_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1594));
   AOI22_X1_50_SVT g79632 (.A0(DPATH_RF_MEMORY_16__21_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__21_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1593));
   AOI22_X1_50_SVT g79633 (.A0(DPATH_RF_MEMORY_9__1_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__1_),
	.B1(n_1399),
	.Q(n_1592));
   AOI22_X1_50_SVT g79634 (.A0(DPATH_RF_MEMORY_13__21_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__21_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1591));
   AO22_X0_50_SVT g79635 (.A0(DPATH_RF_MEMORY_9__21_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__21_),
	.B1(n_1399),
	.Q(n_1590));
   AOI22_X1_50_SVT g79636 (.A0(DPATH_RF_MEMORY_1__12_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__12_),
	.B1(n_1427),
	.Q(n_1589));
   AOI22_X1_50_SVT g79637 (.A0(DPATH_RF_MEMORY_18__12_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__12_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1588));
   AOI22_X1_50_SVT g79638 (.A0(DPATH_RF_MEMORY_21__22_),
	.A1(n_1424),
	.B0(DPATH_RF_MEMORY_22__22_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1587));
   AOI22_X1_50_SVT g79639 (.A0(DPATH_RF_MEMORY_25__20_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__20_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1586));
   AOI22_X1_50_SVT g79640 (.A0(DPATH_RF_MEMORY_24__20_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__20_),
	.B1(n_1445),
	.Q(n_1585));
   AOI22_X1_50_SVT g79641 (.A0(DPATH_RF_MEMORY_29__20_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__20_),
	.B1(n_1378),
	.Q(n_1584));
   AOI22_X1_50_SVT g79642 (.A0(DPATH_RF_MEMORY_28__20_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__20_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1583));
   AOI22_X1_50_SVT g79643 (.A0(DPATH_RF_MEMORY_28__12_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__12_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1582));
   AOI22_X1_50_SVT g79644 (.A0(DPATH_RF_MEMORY_29__12_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__12_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1581));
   AOI22_X1_50_SVT g79645 (.A0(DPATH_RF_MEMORY_9__20_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__20_),
	.B1(n_1399),
	.Q(n_1580));
   AOI22_X1_50_SVT g79646 (.A0(DPATH_RF_MEMORY_24__27_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__27_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1579));
   AOI22_X1_50_SVT g79647 (.A0(DPATH_RF_MEMORY_12__20_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__20_),
	.B1(n_1450),
	.Q(n_1578));
   AOI22_X1_50_SVT g79648 (.A0(DPATH_RF_MEMORY_16__20_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__20_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1577));
   AOI22_X1_50_SVT g79649 (.A0(DPATH_RF_MEMORY_25__12_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__12_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1576));
   AOI22_X1_50_SVT g79650 (.A0(DPATH_RF_MEMORY_1__20_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__20_),
	.B1(n_1434),
	.Q(n_1575));
   AOI22_X1_50_SVT g79651 (.A0(DPATH_RF_MEMORY_5__20_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__20_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1574));
   AOI22_X1_50_SVT g79652 (.A0(DPATH_RF_MEMORY_4__20_),
	.A1(n_1380),
	.B0(DPATH_RF_MEMORY_3__20_),
	.B1(n_1446),
	.Q(n_1573));
   AOI22_X1_50_SVT g79653 (.A0(DPATH_RF_MEMORY_24__12_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__12_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1572));
   AOI22_X1_50_SVT g79654 (.A0(DPATH_RF_MEMORY_17__22_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_31__22_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1571));
   AOI22_X1_50_SVT g79655 (.A0(DPATH_RF_MEMORY_17__11_),
	.A1(n_1414),
	.B0(DPATH_RF_MEMORY_18__11_),
	.B1(FE_OFN57_n_1419),
	.Q(n_1570));
   AOI22_X1_50_SVT g79656 (.A0(DPATH_RF_MEMORY_24__19_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__19_),
	.B1(n_1445),
	.Q(n_1569));
   AOI22_X1_50_SVT g79657 (.A0(DPATH_RF_MEMORY_29__19_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__19_),
	.B1(n_1378),
	.Q(n_1568));
   AOI22_X1_50_SVT g79658 (.A0(DPATH_RF_MEMORY_28__19_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__19_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1567));
   AOI22_X1_50_SVT g79659 (.A0(DPATH_RF_MEMORY_28__22_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__22_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1566));
   AOI22_X1_50_SVT g79660 (.A0(DPATH_RF_MEMORY_25__19_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__19_),
	.B1(n_1389),
	.Q(n_1565));
   AOI22_X1_50_SVT g79661 (.A0(DPATH_RF_MEMORY_20__11_),
	.A1(FE_OFN41_n_1392),
	.B0(DPATH_RF_MEMORY_19__11_),
	.B1(FE_OFN44_n_1396),
	.Q(n_1564));
   AOI22_X1_50_SVT g79662 (.A0(DPATH_RF_MEMORY_12__19_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__19_),
	.B1(n_1450),
	.Q(n_1563));
   AOI22_X1_50_SVT g79663 (.A0(DPATH_RF_MEMORY_13__19_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__19_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1562));
   AOI22_X1_50_SVT g79664 (.A0(DPATH_RF_MEMORY_16__19_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__19_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1561));
   AOI22_X1_50_SVT g79665 (.A0(DPATH_RF_MEMORY_25__22_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__22_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1560));
   AOI22_X1_50_SVT g79666 (.A0(DPATH_RF_MEMORY_5__19_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__19_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1559));
   AOI22_X1_50_SVT g79667 (.A0(DPATH_RF_MEMORY_29__11_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__11_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1558));
   AOI22_X1_50_SVT g79668 (.A0(DPATH_RF_MEMORY_8__19_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__19_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1557));
   AOI22_X1_50_SVT g79669 (.A0(DPATH_RF_MEMORY_4__19_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__19_),
	.B1(n_1446),
	.Q(n_1556));
   AOI22_X1_50_SVT g79670 (.A0(DPATH_RF_MEMORY_8__31_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__31_),
	.B1(n_1403),
	.Q(n_1555));
   AOI22_X1_50_SVT g79671 (.A0(DPATH_RF_MEMORY_20__18_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_31__18_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1554));
   AOI22_X1_50_SVT g79672 (.A0(DPATH_RF_MEMORY_13__27_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__27_),
	.B1(n_1412),
	.Q(n_1553));
   AOI22_X1_50_SVT g79673 (.A0(DPATH_RF_MEMORY_25__11_),
	.A1(FE_OFN45_n_1397),
	.B0(DPATH_RF_MEMORY_26__11_),
	.B1(FE_OFN53_n_1409),
	.Q(n_1552));
   AOI22_X1_50_SVT g79674 (.A0(DPATH_RF_MEMORY_13__2_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__2_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1551));
   AOI22_X1_50_SVT g79675 (.A0(DPATH_RF_MEMORY_28__11_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__11_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1550));
   AOI22_X1_50_SVT g79676 (.A0(DPATH_RF_MEMORY_13__18_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__18_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1549));
   AOI22_X1_50_SVT g79677 (.A0(DPATH_RF_MEMORY_12__18_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__18_),
	.B1(n_1450),
	.Q(n_1548));
   AOI22_X1_50_SVT g79678 (.A0(DPATH_RF_MEMORY_16__18_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__18_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1547));
   AOI22_X1_50_SVT g79679 (.A0(DPATH_RF_MEMORY_9__18_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__18_),
	.B1(n_1399),
	.Q(n_1546));
   AOI22_X1_50_SVT g79680 (.A0(DPATH_RF_MEMORY_24__11_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__11_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1545));
   AO22_X0_50_SVT g79681 (.A0(DPATH_RF_MEMORY_24__22_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__22_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1544));
   AOI22_X1_50_SVT g79682 (.A0(DPATH_RF_MEMORY_24__18_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__18_),
	.B1(n_1445),
	.Q(n_1543));
   AOI22_X1_50_SVT g79683 (.A0(DPATH_RF_MEMORY_28__18_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__18_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1542));
   AOI22_X1_50_SVT g79684 (.A0(DPATH_RF_MEMORY_16__27_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__27_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1541));
   AOI22_X1_50_SVT g79685 (.A0(DPATH_RF_MEMORY_1__18_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__18_),
	.B1(n_1434),
	.Q(n_1540));
   AOI22_X1_50_SVT g79686 (.A0(DPATH_RF_MEMORY_8__18_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__18_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1539));
   AOI22_X1_50_SVT g79687 (.A0(DPATH_RF_MEMORY_16__29_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__29_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1538));
   AO22_X0_50_SVT g79688 (.A0(DPATH_RF_MEMORY_5__18_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__18_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1537));
   AOI22_X1_50_SVT g79689 (.A0(DPATH_RF_MEMORY_5__11_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__11_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1536));
   AOI22_X1_50_SVT g79690 (.A0(DPATH_RF_MEMORY_1__17_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__17_),
	.B1(n_1434),
	.Q(n_1535));
   AOI22_X1_50_SVT g79691 (.A0(DPATH_RF_MEMORY_4__21_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__21_),
	.B1(n_1420),
	.Q(n_1534));
   AOI22_X1_50_SVT g79692 (.A0(DPATH_RF_MEMORY_5__17_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__17_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1533));
   AOI22_X1_50_SVT g79693 (.A0(DPATH_RF_MEMORY_1__11_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__11_),
	.B1(n_1427),
	.Q(n_1532));
   AOI22_X1_50_SVT g79694 (.A0(DPATH_RF_MEMORY_8__17_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__17_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1531));
   AOI22_X1_50_SVT g79695 (.A0(DPATH_RF_MEMORY_4__17_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__17_),
	.B1(n_1446),
	.Q(n_1530));
   AOI22_X1_50_SVT g79696 (.A0(DPATH_RF_MEMORY_9__11_),
	.A1(FE_PDN1443_FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__11_),
	.B1(n_1417),
	.Q(n_1529));
   AOI22_X1_50_SVT g79697 (.A0(DPATH_RF_MEMORY_1__27_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__27_),
	.B1(n_1427),
	.Q(n_1528));
   AOI22_X1_50_SVT g79698 (.A0(DPATH_RF_MEMORY_25__17_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__17_),
	.B1(n_1389),
	.Q(n_1527));
   AOI22_X1_50_SVT g79699 (.A0(DPATH_RF_MEMORY_29__17_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__17_),
	.B1(n_1378),
	.Q(n_1526));
   AOI22_X1_50_SVT g79700 (.A0(DPATH_RF_MEMORY_28__17_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__17_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1525));
   AOI22_X1_50_SVT g79701 (.A0(DPATH_RF_MEMORY_13__11_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__11_),
	.B1(n_1412),
	.Q(n_1524));
   AOI22_X1_50_SVT g79702 (.A0(DPATH_RF_MEMORY_17__17_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__17_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1523));
   AOI22_X1_50_SVT g79703 (.A0(DPATH_RF_MEMORY_21__17_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__17_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1522));
   AOI22_X1_50_SVT g79704 (.A0(DPATH_RF_MEMORY_12__11_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__11_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1521));
   AOI22_X1_50_SVT g79705 (.A0(DPATH_RF_MEMORY_9__17_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__17_),
	.B1(n_1399),
	.Q(n_1520));
   AOI22_X1_50_SVT g79706 (.A0(DPATH_RF_MEMORY_16__17_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__17_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1519));
   AOI22_X1_50_SVT g79707 (.A0(DPATH_RF_MEMORY_1__21_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__21_),
	.B1(n_1427),
	.Q(n_1518));
   AO22_X0_50_SVT g79708 (.A0(DPATH_RF_MEMORY_13__17_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__17_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1517));
   AOI22_X1_50_SVT g79709 (.A0(DPATH_RF_MEMORY_16__11_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__11_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1516));
   AOI22_X1_50_SVT g79710 (.A0(DPATH_RF_MEMORY_5__21_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__21_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1515));
   AOI22_X1_50_SVT g79711 (.A0(DPATH_RF_MEMORY_8__21_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__21_),
	.B1(n_1403),
	.Q(n_1514));
   AOI22_X1_50_SVT g79712 (.A0(DPATH_RF_MEMORY_5__16_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__16_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1513));
   AOI22_X1_50_SVT g79713 (.A0(DPATH_RF_MEMORY_5__10_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__10_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1512));
   AOI22_X1_50_SVT g79714 (.A0(DPATH_RF_MEMORY_4__16_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__16_),
	.B1(n_1446),
	.Q(n_1511));
   AOI22_X1_50_SVT g79715 (.A0(DPATH_RF_MEMORY_8__8_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__8_),
	.B1(n_1403),
	.Q(n_1510));
   AOI22_X1_50_SVT g79716 (.A0(DPATH_RF_MEMORY_4__27_),
	.A1(FE_OFN58_n_1422),
	.B0(DPATH_RF_MEMORY_3__27_),
	.B1(n_1420),
	.Q(n_1509));
   AOI22_X1_50_SVT g79717 (.A0(DPATH_RF_MEMORY_8__16_),
	.A1(n_1444),
	.B0(DPATH_RF_MEMORY_7__16_),
	.B1(FE_OFN69_n_1443),
	.Q(n_1508));
   AOI22_X1_50_SVT g79718 (.A0(DPATH_RF_MEMORY_1__16_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__16_),
	.B1(n_1434),
	.Q(n_1507));
   AOI22_X1_50_SVT g79719 (.A0(DPATH_RF_MEMORY_29__16_),
	.A1(n_1406),
	.B0(DPATH_RF_MEMORY_30__16_),
	.B1(n_1378),
	.Q(n_1506));
   AOI22_X1_50_SVT g79720 (.A0(DPATH_RF_MEMORY_25__16_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__16_),
	.B1(FE_OFN38_n_1389),
	.Q(n_1505));
   AOI22_X1_50_SVT g79721 (.A0(DPATH_RF_MEMORY_24__16_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__16_),
	.B1(n_1445),
	.Q(n_1504));
   AOI22_X1_50_SVT g79722 (.A0(DPATH_RF_MEMORY_8__10_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__10_),
	.B1(n_1403),
	.Q(n_1503));
   AOI22_X1_50_SVT g79723 (.A0(DPATH_RF_MEMORY_17__16_),
	.A1(FE_OFN26_n_1371),
	.B0(DPATH_RF_MEMORY_31__16_),
	.B1(FE_OFN36_n_1386),
	.Q(n_1502));
   AOI22_X1_50_SVT g79724 (.A0(DPATH_RF_MEMORY_21__16_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__16_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1501));
   AO22_X0_50_SVT g79725 (.A0(DPATH_RF_MEMORY_1__10_),
	.A1(FE_OFN28_n_1376),
	.B0(DPATH_RF_MEMORY_2__10_),
	.B1(n_1427),
	.Q(n_1500));
   AOI22_X1_50_SVT g79726 (.A0(DPATH_RF_MEMORY_9__16_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__16_),
	.B1(n_1399),
	.Q(n_1499));
   AOI22_X1_50_SVT g79727 (.A0(DPATH_RF_MEMORY_12__16_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__16_),
	.B1(n_1450),
	.Q(n_1498));
   AO22_X0_50_SVT g79728 (.A0(DPATH_RF_MEMORY_16__16_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__16_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1497));
   AOI22_X1_50_SVT g79729 (.A0(DPATH_RF_MEMORY_5__27_),
	.A1(n_1410),
	.B0(DPATH_RF_MEMORY_6__27_),
	.B1(FE_OFN59_n_1423),
	.Q(n_1496));
   AOI22_X1_50_SVT g79730 (.A0(DPATH_RF_MEMORY_16__15_),
	.A1(n_1447),
	.B0(DPATH_RF_MEMORY_15__15_),
	.B1(FE_OFN72_n_1448),
	.Q(n_1495));
   AOI22_X1_50_SVT g79731 (.A0(DPATH_RF_MEMORY_12__11_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__11_),
	.B1(n_1450),
	.Q(n_1494));
   AOI22_X1_50_SVT g79732 (.A0(DPATH_RF_MEMORY_9__15_),
	.A1(n_1430),
	.B0(DPATH_RF_MEMORY_10__15_),
	.B1(n_1399),
	.Q(n_1493));
   AOI22_X1_50_SVT g79733 (.A0(DPATH_RF_MEMORY_13__15_),
	.A1(FE_OFN73_n_1449),
	.B0(DPATH_RF_MEMORY_14__15_),
	.B1(FE_OFN48_n_1401),
	.Q(n_1492));
   AOI22_X1_50_SVT g79734 (.A0(DPATH_RF_MEMORY_12__15_),
	.A1(FE_OFN47_n_1400),
	.B0(DPATH_RF_MEMORY_11__15_),
	.B1(n_1450),
	.Q(n_1491));
   AOI22_X1_50_SVT g79735 (.A0(DPATH_RF_MEMORY_9__29_),
	.A1(FE_OFN34_n_1383),
	.B0(DPATH_RF_MEMORY_10__29_),
	.B1(n_1417),
	.Q(n_1490));
   AOI22_X1_50_SVT g79736 (.A0(DPATH_RF_MEMORY_21__10_),
	.A1(n_1425),
	.B0(DPATH_RF_MEMORY_22__10_),
	.B1(FE_OFN25_n_1331),
	.Q(n_1489));
   AOI22_X1_50_SVT g79737 (.A0(DPATH_RF_MEMORY_4__15_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__15_),
	.B1(n_1446),
	.Q(n_1488));
   AOI22_X1_50_SVT g79738 (.A0(DPATH_RF_MEMORY_5__15_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__15_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1487));
   AOI22_X1_50_SVT g79739 (.A0(DPATH_RF_MEMORY_28__21_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__21_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1486));
   AOI22_X1_50_SVT g79740 (.A0(DPATH_RF_MEMORY_1__15_),
	.A1(n_1372),
	.B0(DPATH_RF_MEMORY_2__15_),
	.B1(n_1434),
	.Q(n_1485));
   AOI22_X1_50_SVT g79741 (.A0(DPATH_RF_MEMORY_13__10_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__10_),
	.B1(n_1412),
	.Q(n_1484));
   AOI22_X1_50_SVT g79742 (.A0(DPATH_RF_MEMORY_29__21_),
	.A1(FE_OFN39_n_1390),
	.B0(DPATH_RF_MEMORY_30__21_),
	.B1(FE_OFN29_n_1377),
	.Q(n_1483));
   AOI22_X1_50_SVT g79743 (.A0(DPATH_RF_MEMORY_20__15_),
	.A1(FE_OFN52_n_1408),
	.B0(DPATH_RF_MEMORY_19__15_),
	.B1(FE_OFN66_n_1440),
	.Q(n_1482));
   AOI22_X1_50_SVT g79744 (.A0(DPATH_RF_MEMORY_8__27_),
	.A1(FE_OFN27_n_1374),
	.B0(DPATH_RF_MEMORY_7__27_),
	.B1(n_1403),
	.Q(n_1481));
   AOI22_X1_50_SVT g79745 (.A0(DPATH_RF_MEMORY_13__29_),
	.A1(FE_OFN42_n_1393),
	.B0(DPATH_RF_MEMORY_14__29_),
	.B1(n_1412),
	.Q(n_1480));
   AOI22_X1_50_SVT g79746 (.A0(DPATH_RF_MEMORY_12__10_),
	.A1(n_1421),
	.B0(DPATH_RF_MEMORY_11__10_),
	.B1(FE_OFN40_n_1391),
	.Q(n_1479));
   AOI22_X1_50_SVT g79747 (.A0(DPATH_RF_MEMORY_21__15_),
	.A1(FE_OFN64_n_1436),
	.B0(DPATH_RF_MEMORY_22__15_),
	.B1(FE_OFN65_n_1438),
	.Q(n_1478));
   AOI22_X1_50_SVT g79748 (.A0(DPATH_RF_MEMORY_24__21_),
	.A1(FE_OFN46_n_1398),
	.B0(DPATH_RF_MEMORY_23__21_),
	.B1(FE_OFN33_n_1381),
	.Q(n_1477));
   AOI22_X1_50_SVT g79749 (.A0(DPATH_RF_MEMORY_25__15_),
	.A1(FE_OFN68_n_1442),
	.B0(DPATH_RF_MEMORY_26__15_),
	.B1(n_1389),
	.Q(n_1476));
   AOI22_X1_50_SVT g79750 (.A0(DPATH_RF_MEMORY_28__6_),
	.A1(FE_OFN54_n_1411),
	.B0(DPATH_RF_MEMORY_27__6_),
	.B1(FE_OFN55_n_1413),
	.Q(n_1475));
   AOI22_X1_50_SVT g79751 (.A0(DPATH_RF_MEMORY_24__15_),
	.A1(n_1405),
	.B0(DPATH_RF_MEMORY_23__15_),
	.B1(n_1445),
	.Q(n_1474));
   AO22_X0_50_SVT g79752 (.A0(DPATH_RF_MEMORY_28__15_),
	.A1(FE_OFN67_n_1441),
	.B0(DPATH_RF_MEMORY_27__15_),
	.B1(FE_OFN31_n_1379),
	.Q(n_1473));
   AOI22_X1_50_SVT g79753 (.A0(DPATH_RF_MEMORY_16__10_),
	.A1(FE_OFN43_n_1395),
	.B0(DPATH_RF_MEMORY_15__10_),
	.B1(FE_OFN62_n_1429),
	.Q(n_1472));
   AOI22_X1_50_SVT g79754 (.A0(DPATH_RF_MEMORY_5__14_),
	.A1(n_1387),
	.B0(DPATH_RF_MEMORY_6__14_),
	.B1(FE_OFN49_n_1404),
	.Q(n_1471));
   AOI22_X1_50_SVT g79755 (.A0(DPATH_RF_MEMORY_18__10_),
	.A1(FE_OFN57_n_1419),
	.B0(DPATH_RF_MEMORY_31__10_),
	.B1(FE_OFN35_n_1385),
	.Q(n_1470));
   AOI22_X1_50_SVT g79756 (.A0(DPATH_RF_MEMORY_4__14_),
	.A1(FE_OFN32_n_1380),
	.B0(DPATH_RF_MEMORY_3__14_),
	.B1(n_1446),
	.Q(n_1469));
   CLKNAND2_X2_50_SVT g79758 (.A(DPATH_RF_MEMORY_20__2_),
	.B(n_1408),
	.Q(n_1466));
   CLKNAND2_X2_50_SVT g79759 (.A(DPATH_RF_MEMORY_31__11_),
	.B(FE_OFN36_n_1386),
	.Q(n_1465));
   CLKNAND2_X2_50_SVT g79760 (.A(DPATH_RF_MEMORY_21__5_),
	.B(n_1436),
	.Q(n_1464));
   CLKNAND2_X2_50_SVT g79761 (.A(DPATH_RF_MEMORY_31__1_),
	.B(n_1386),
	.Q(n_1463));
   NAND2T_X1_50_SVT g79762 (.A(DPATH_RF_MEMORY_17__19_),
	.B(n_1414),
	.Q(n_1462));
   NAND2T_X1_50_SVT g79763 (.A(DPATH_RF_MEMORY_18__18_),
	.B(FE_OFN57_n_1419),
	.Q(n_1461));
   NAND2_X0_50_SVT g79764 (.A(n_1352),
	.B(n_1451),
	.Q(n_1468));
   NAND2T_X1_50_SVT g79765 (.A(DPATH_RF_MEMORY_20__5_),
	.B(FE_OFN41_n_1392),
	.Q(n_1460));
   CLKNAND2_X2_50_SVT g79766 (.A(DPATH_RF_MEMORY_21__9_),
	.B(n_1436),
	.Q(n_1459));
   NAND2T_X1_50_SVT g79767 (.A(DPATH_RF_MEMORY_21__17_),
	.B(n_1424),
	.Q(n_1458));
   CLKNAND2_X2_50_SVT g79768 (.A(DPATH_RF_MEMORY_17__18_),
	.B(FE_OFN26_n_1371),
	.Q(n_1457));
   CLKNAND2_X2_50_SVT g79769 (.A(DPATH_RF_MEMORY_19__4_),
	.B(FE_OFN66_n_1440),
	.Q(n_1456));
   CLKNAND2_X2_50_SVT g79770 (.A(DPATH_RF_MEMORY_20__25_),
	.B(FE_OFN52_n_1408),
	.Q(n_1455));
   CLKNAND2_X2_50_SVT g79771 (.A(DPATH_RF_MEMORY_31__13_),
	.B(n_1386),
	.Q(n_1454));
   CLKNAND2_X2_50_SVT g79772 (.A(DPATH_RF_MEMORY_21__24_),
	.B(FE_OFN64_n_1436),
	.Q(n_1453));
   NAND2T_X1_50_SVT g79773 (.A(DPATH_RF_MEMORY_20__25_),
	.B(FE_OFN41_n_1392),
	.Q(n_1452));
   INV_X4_50_SVT g79777 (.A(n_1433),
	.Q(n_1434));
   CLKINV_X6_50_SVT g79783 (.A(n_1416),
	.Q(n_1417));
   NOR2_X0_50_SVT g79785 (.A(INSTR[2]),
	.B(MEMWRITE),
	.Q(n_1451));
   AND2_X4_50_SVT g79786 (.A(n_1360),
	.B(n_1349),
	.Q(n_1450));
   INV_A_NOR2_X0_50_SVT g79787 (.AN(n_1329),
	.B(n_1345),
	.Q(n_1449));
   INV_A_NOR2_X0_50_SVT g79788 (.AN(n_1360),
	.B(n_1345),
	.Q(n_1448));
   NOR2P3_X6_50_SVT g79789 (.A(n_1361),
	.B(n_1337),
	.Q(n_1447));
   AND2_X4_50_SVT g79790 (.A(n_1326),
	.B(n_1349),
	.Q(n_1446));
   NOR2P3T_X4_50_SVT g79791 (.A(n_1362),
	.B(n_1345),
	.Q(n_1445));
   AND2_X4_50_SVT g79792 (.A(n_1329),
	.B(n_1338),
	.Q(n_1444));
   INV_A_NOR2_X0_50_SVT g79793 (.AN(n_1326),
	.B(n_1345),
	.Q(n_1443));
   NOR2_X0_50_SVT g79794 (.A(n_1350),
	.B(n_1367),
	.Q(n_1442));
   NOR2_X0_50_SVT g79795 (.A(n_1367),
	.B(n_1346),
	.Q(n_1441));
   NOR2P3_X2_50_SVT g79796 (.A(n_1350),
	.B(n_1362),
	.Q(n_1440));
   NOR2_X0_50_SVT g79797 (.A(n_1362),
	.B(n_1346),
	.Q(n_1438));
   NOR2P3_X2_50_SVT g79798 (.A(n_1345),
	.B(n_1361),
	.Q(n_1436));
   NAND2_X0_50_SVT g79799 (.A(n_1338),
	.B(n_1326),
	.Q(n_1433));
   NOR2_X0_50_SVT g79800 (.A(n_1362),
	.B(n_1337),
	.Q(n_1432));
   AND2_X4_50_SVT g79801 (.A(n_1329),
	.B(n_1349),
	.Q(n_1430));
   INV_A_NOR2_X0_50_SVT g79802 (.AN(n_1363),
	.B(n_1351),
	.Q(n_1429));
   CLKAND2_X4_50_SVT g79803 (.A(n_1328),
	.B(n_1339),
	.Q(n_1427));
   NOR2P3_X2_50_SVT g79804 (.A(n_1334),
	.B(n_1358),
	.Q(n_1425));
   AND2_X0_50_SVT g79805 (.A(n_1363),
	.B(n_1339),
	.Q(n_1423));
   AND2_X0_50_SVT g79806 (.A(n_1327),
	.B(n_1339),
	.Q(n_1422));
   AND2_X4_50_SVT g79807 (.A(n_1327),
	.B(n_1348),
	.Q(n_1421));
   CLKAND2_X4_50_SVT g79808 (.A(n_1328),
	.B(n_1335),
	.Q(n_1420));
   INV_A_NAND2_X0_50_SVT g79809 (.AN(n_1364),
	.B(n_1339),
	.Q(n_1419));
   NAND2_X1_50_SVT g79810 (.A(n_1348),
	.B(n_1328),
	.Q(n_1416));
   NOR2P3_X2_50_SVT g79811 (.A(n_1334),
	.B(n_1357),
	.Q(n_1415));
   NOR2_X0_50_SVT g79812 (.A(n_1364),
	.B(n_1351),
	.Q(n_1413));
   AND2_X4_50_SVT g79813 (.A(n_1363),
	.B(n_1348),
	.Q(n_1412));
   NOR2_X0_50_SVT g79814 (.A(n_1358),
	.B(n_1347),
	.Q(n_1411));
   AND2_X4_50_SVT g79815 (.A(n_1327),
	.B(n_1335),
	.Q(n_1410));
   NOR2_X0_50_SVT g79816 (.A(n_1364),
	.B(n_1347),
	.Q(n_1409));
   NOR2P3_X2_50_SVT g79828 (.A(n_1346),
	.B(n_1361),
	.Q(n_1408));
   NOR2P3T_X4_50_SVT g79829 (.A(n_1345),
	.B(n_1367),
	.Q(n_1406));
   NOR2P3T_X4_50_SVT g79830 (.A(n_1337),
	.B(n_1367),
	.Q(n_1405));
   INV_A_NOR2_X0_50_SVT g79831 (.AN(n_1326),
	.B(n_1346),
	.Q(n_1404));
   CLKAND2_X4_50_SVT g79832 (.A(n_1363),
	.B(n_1335),
	.Q(n_1403));
   INV_A_NOR2_X0_50_SVT g79833 (.AN(n_1360),
	.B(n_1346),
	.Q(n_1401));
   INV_A_NOR2_X0_50_SVT g79834 (.AN(n_1329),
	.B(n_1346),
	.Q(n_1400));
   AND2_X4_50_SVT g79835 (.A(n_1360),
	.B(n_1338),
	.Q(n_1399));
   NOR2_X0_50_SVT g79836 (.A(n_1357),
	.B(n_1347),
	.Q(n_1398));
   NOR2_X0_50_SVT g79837 (.A(n_1357),
	.B(n_1351),
	.Q(n_1397));
   NOR2_X0_50_SVT g79838 (.A(n_1364),
	.B(n_1334),
	.Q(n_1396));
   INV_A_NOR2_X1_50_SVT g79839 (.AN(n_1339),
	.B(n_1357),
	.Q(n_1395));
   INV_A_NOR2_X0_50_SVT g79840 (.AN(n_1327),
	.B(n_1351),
	.Q(n_1393));
   INV_A_NOR2_X1_50_SVT g79841 (.AN(n_1339),
	.B(n_1358),
	.Q(n_1392));
   INV_A_NOR2_X0_50_SVT g79842 (.AN(n_1328),
	.B(n_1351),
	.Q(n_1391));
   NOR2_X0_50_SVT g79843 (.A(n_1351),
	.B(n_1358),
	.Q(n_1390));
   NOR2P3T_X2_50_SVT g79844 (.A(n_1366),
	.B(n_1337),
	.Q(n_1389));
   NOR2P3T_X4_50_SVT g79846 (.A(n_1345),
	.B(n_1368),
	.Q(n_1387));
   NOR2P3_X2_50_SVT g79847 (.A(n_1366),
	.B(n_1345),
	.Q(n_1386));
   NOR2_X0_50_SVT g79848 (.A(n_1365),
	.B(n_1351),
	.Q(n_1385));
   NOR2_X0_50_SVT g79849 (.A(n_1351),
	.B(n_1369),
	.Q(n_1383));
   NOR2_X0_50_SVT g79850 (.A(n_1365),
	.B(n_1334),
	.Q(n_1381));
   NOR2P3_X2_50_SVT g79851 (.A(n_1346),
	.B(n_1368),
	.Q(n_1380));
   NOR2_X0_50_SVT g79852 (.A(n_1366),
	.B(n_1350),
	.Q(n_1379));
   NOR2P3T_X4_50_SVT g79853 (.A(n_1366),
	.B(n_1346),
	.Q(n_1378));
   NOR2_X0_50_SVT g79854 (.A(n_1365),
	.B(n_1347),
	.Q(n_1377));
   NOR2_X0_50_SVT g79855 (.A(n_1369),
	.B(n_1334),
	.Q(n_1376));
   NOR2_X0_50_SVT g79856 (.A(n_1369),
	.B(n_1347),
	.Q(n_1374));
   NOR2P3_X2_50_SVT g79858 (.A(n_1350),
	.B(n_1361),
	.Q(n_1371));
   INV_A_NAND2_X0_50_SVT g79861 (.AN(INSTR[24]),
	.B(n_1343),
	.Q(n_1369));
   INV_A_NAND2_X0_50_SVT g79862 (.AN(INSTR[19]),
	.B(n_1353),
	.Q(n_1368));
   NAND2_X0_50_SVT g79864 (.A(INSTR[19]),
	.B(n_1354),
	.Q(n_1367));
   INV_A_NAND2_X0_50_SVT g79865 (.AN(n_1341),
	.B(INSTR[19]),
	.Q(n_1366));
   INV_A_NAND2_X0_50_SVT g79867 (.AN(n_1355),
	.B(INSTR[24]),
	.Q(n_1365));
   NAND2_X0_50_SVT g79868 (.A(INSTR[24]),
	.B(n_1344),
	.Q(n_1364));
   NOR2_X0_50_SVT g79869 (.A(INSTR[24]),
	.B(n_1355),
	.Q(n_1363));
   NAND2_X0_50_SVT g79871 (.A(INSTR[19]),
	.B(n_1340),
	.Q(n_1362));
   NAND2_X0_50_SVT g79872 (.A(INSTR[19]),
	.B(n_1353),
	.Q(n_1361));
   NOR2_X0_50_SVT g79873 (.A(INSTR[19]),
	.B(n_1341),
	.Q(n_1360));
   INV_A_OAI21_X0_50_SVT g79876 (.A0(n_3),
	.A1N(INSTR[16]),
	.B0(n_1336),
	.Q(DPATH_n_5214));
   INV_A_OAI21_X0_50_SVT g79877 (.A0(n_3),
	.A1N(INSTR[13]),
	.B0(n_1336),
	.Q(DPATH_n_5217));
   INV_A_OAI21_X0_50_SVT g79878 (.A0(n_3),
	.A1N(INSTR[12]),
	.B0(n_1336),
	.Q(DPATH_n_5218));
   INV_A_OAI21_X0_50_SVT g79879 (.A0(n_3),
	.A1N(INSTR[14]),
	.B0(n_1336),
	.Q(DPATH_n_5216));
   INV_A_OAI21_X0_50_SVT g79880 (.A0(n_3),
	.A1N(INSTR[18]),
	.B0(n_1336),
	.Q(DPATH_n_5212));
   INV_A_OAI21_X0_50_SVT g79881 (.A0(n_3),
	.A1N(INSTR[15]),
	.B0(n_1336),
	.Q(DPATH_n_5215));
   INV_A_OAI21_X0_50_SVT g79882 (.A0(n_3),
	.A1N(INSTR[17]),
	.B0(n_1336),
	.Q(DPATH_n_5213));
   INV_A_OAI21_X0_50_SVT g79883 (.A0(n_3),
	.A1N(INSTR[19]),
	.B0(n_1336),
	.Q(DPATH_n_5211));
   INV_A_NOR3_X2_50_SVT g79884 (.AN(INSTR[5]),
	.B(INSTR[6]),
	.C(INSTR[4]),
	.Q(MEMWRITE));
   NAND2_X0_50_SVT g79885 (.A(INSTR[24]),
	.B(n_1342),
	.Q(n_1358));
   NAND2_X0_50_SVT g79886 (.A(INSTR[24]),
	.B(n_1343),
	.Q(n_1357));
   CLKNAND2_X4_50_SVT g79888 (.A(n_1352),
	.B(n_2708),
	.Q(n_1356));
   NAND2_X0_50_SVT g79892 (.A(INSTR[21]),
	.B(INSTR[22]),
	.Q(n_1355));
   INV_A_NOR2_X0_50_SVT g79893 (.AN(INSTR[18]),
	.B(INSTR[16]),
	.Q(n_1354));
   NAND2_X0_50_SVT g79894 (.A(INSTR[4]),
	.B(INSTR[5]),
	.Q(n_2708));
   NOR2_X0_50_SVT g79895 (.A(INSTR[16]),
	.B(INSTR[18]),
	.Q(n_1353));
   NOR2_X0_50_SVT g79896 (.A(INSTR[2]),
	.B(INSTR[6]),
	.Q(n_1352));
   NAND2_X1_50_SVT g79897 (.A(INSTR[23]),
	.B(INSTR[20]),
	.Q(n_1351));
   INV_A_NAND2_X0_50_SVT g79898 (.AN(INSTR[17]),
	.B(INSTR[15]),
	.Q(n_1350));
   INV_A_NOR2_X0_50_SVT g79899 (.AN(INSTR[23]),
	.B(INSTR[20]),
	.Q(n_1348));
   INV_A_NAND2_X1_50_SVT g79900 (.AN(INSTR[15]),
	.B(INSTR[17]),
	.Q(n_1346));
   NAND2_X1_50_SVT g79901 (.A(INSTR[17]),
	.B(INSTR[15]),
	.Q(n_1345));
   NAND2_X0_50_SVT g79907 (.A(INSTR[6]),
	.B(n_3),
	.Q(n_2706));
   INV_A_NOR2_X0_50_SVT g79908 (.AN(INSTR[21]),
	.B(INSTR[22]),
	.Q(n_1344));
   NOR2_X0_50_SVT g79909 (.A(INSTR[21]),
	.B(INSTR[22]),
	.Q(n_1343));
   INV_A_NOR2_X0_50_SVT g79910 (.AN(INSTR[22]),
	.B(INSTR[21]),
	.Q(n_1342));
   NAND2_X0_50_SVT g79911 (.A(INSTR[16]),
	.B(INSTR[18]),
	.Q(n_1341));
   INV_A_NOR2_X0_50_SVT g79912 (.AN(INSTR[16]),
	.B(INSTR[18]),
	.Q(n_1340));
   NOR2_X0_50_SVT g79913 (.A(INSTR[20]),
	.B(INSTR[23]),
	.Q(n_1339));
   NOR2_X0_50_SVT g79914 (.A(INSTR[15]),
	.B(INSTR[17]),
	.Q(n_1338));
   NAND2_X0_50_SVT g79915 (.A(INSTR[31]),
	.B(n_3),
	.Q(n_1336));
   INV_A_NOR2_X0_50_SVT g79916 (.AN(INSTR[20]),
	.B(INSTR[23]),
	.Q(n_1335));
   INV_X2_50_SVT g79917 (.A(INSTR[2]),
	.Q(n_3));
   INV_A_NAND2_X0_50_SVT g2 (.AN(n_1368),
	.B(n_1349),
	.Q(n_1332));
   INV_A_NOR2_X0_50_SVT g79918 (.AN(n_1339),
	.B(n_1365),
	.Q(n_1331));
   INV_A_NAND2_X2_50_SVT g79919 (.AN(n_1356),
	.B(INSTR[31]),
	.Q(n_1330));
   INV_A_NOR2_X2_50_SVT g79920 (.AN(n_1354),
	.B(INSTR[19]),
	.Q(n_1329));
   INV_A_NOR2_X2_50_SVT g79921 (.AN(n_1344),
	.B(INSTR[24]),
	.Q(n_1328));
   INV_A_NOR2_X2_50_SVT g79922 (.AN(n_1342),
	.B(INSTR[24]),
	.Q(n_1327));
   INV_A_NOR2_X2_50_SVT g79923 (.AN(n_1340),
	.B(INSTR[19]),
	.Q(n_1326));
   XOR3_X2_50_SVT g28748 (.A(DPATH_n_2758),
	.B(DPATH_n_2796),
	.C(n_1325),
	.Q(ALURSLT[31]));
   FA1_X1_50_SVT g28749 (.A(DPATH_n_2797),
	.B(DPATH_n_2759),
	.CI(n_1324),
	.CO(n_1325),
	.S(ALURSLT[30]));
   FA1_X1_50_SVT g28750 (.A(DPATH_n_2798),
	.B(DPATH_n_2760),
	.CI(n_1323),
	.CO(n_1324),
	.S(ALURSLT[29]));
   FA1_X1_50_SVT g28751 (.A(DPATH_n_2799),
	.B(DPATH_n_2761),
	.CI(n_1322),
	.CO(n_1323),
	.S(ALURSLT[28]));
   FA1_X1_50_SVT g28752 (.A(DPATH_n_2800),
	.B(DPATH_n_2762),
	.CI(n_1321),
	.CO(n_1322),
	.S(ALURSLT[27]));
   FA1_X1_50_SVT g28753 (.A(DPATH_n_2801),
	.B(DPATH_n_2763),
	.CI(n_1320),
	.CO(n_1321),
	.S(ALURSLT[26]));
   FA1_X1_50_SVT g28754 (.A(DPATH_n_2802),
	.B(DPATH_n_2764),
	.CI(n_1319),
	.CO(n_1320),
	.S(ALURSLT[25]));
   FA1_X1_50_SVT g28755 (.A(DPATH_n_2803),
	.B(DPATH_n_2765),
	.CI(n_1318),
	.CO(n_1319),
	.S(ALURSLT[24]));
   FA1_X1_50_SVT g28756 (.A(DPATH_n_2804),
	.B(DPATH_n_2766),
	.CI(n_1317),
	.CO(n_1318),
	.S(ALURSLT[23]));
   FA1_X1_50_SVT g28757 (.A(DPATH_n_2805),
	.B(DPATH_n_2767),
	.CI(n_1316),
	.CO(n_1317),
	.S(ALURSLT[22]));
   FA1_X1_50_SVT g28758 (.A(DPATH_n_2806),
	.B(DPATH_n_2768),
	.CI(n_1315),
	.CO(n_1316),
	.S(ALURSLT[21]));
   FA1_X1_50_SVT g28759 (.A(DPATH_n_2807),
	.B(DPATH_n_2769),
	.CI(n_1314),
	.CO(n_1315),
	.S(ALURSLT[20]));
   FA1_X1_50_SVT g28760 (.A(DPATH_n_2808),
	.B(DPATH_n_2770),
	.CI(n_1313),
	.CO(n_1314),
	.S(ALURSLT[19]));
   FA1_X1_50_SVT g28761 (.A(DPATH_n_2809),
	.B(DPATH_n_2771),
	.CI(n_1312),
	.CO(n_1313),
	.S(ALURSLT[18]));
   FA1_X1_50_SVT g28762 (.A(DPATH_n_2810),
	.B(DPATH_n_2772),
	.CI(n_1311),
	.CO(n_1312),
	.S(ALURSLT[17]));
   FA1_X1_50_SVT g28763 (.A(DPATH_n_2811),
	.B(DPATH_n_2773),
	.CI(n_1310),
	.CO(n_1311),
	.S(ALURSLT[16]));
   FA1_X1_50_SVT g28764 (.A(DPATH_n_2812),
	.B(DPATH_n_2774),
	.CI(n_1309),
	.CO(n_1310),
	.S(ALURSLT[15]));
   FA1_X1_50_SVT g28765 (.A(DPATH_n_2813),
	.B(DPATH_n_2775),
	.CI(n_1308),
	.CO(n_1309),
	.S(ALURSLT[14]));
   FA1_X1_50_SVT g28766 (.A(DPATH_n_2814),
	.B(DPATH_n_2776),
	.CI(n_1307),
	.CO(n_1308),
	.S(ALURSLT[13]));
   FA1_X1_50_SVT g28767 (.A(DPATH_n_2815),
	.B(DPATH_n_2777),
	.CI(n_1306),
	.CO(n_1307),
	.S(ALURSLT[12]));
   FA1_X1_50_SVT g28768 (.A(DPATH_n_2816),
	.B(DPATH_n_2778),
	.CI(n_1305),
	.CO(n_1306),
	.S(ALURSLT[11]));
   FA1_X1_50_SVT g28769 (.A(DPATH_n_2817),
	.B(DPATH_n_2779),
	.CI(n_1304),
	.CO(n_1305),
	.S(ALURSLT[10]));
   FA1_X1_50_SVT g28770 (.A(DPATH_n_2818),
	.B(DPATH_n_2780),
	.CI(n_1303),
	.CO(n_1304),
	.S(ALURSLT[9]));
   FA1_X1_50_SVT g28771 (.A(DPATH_n_2819),
	.B(DPATH_n_2781),
	.CI(n_1302),
	.CO(n_1303),
	.S(ALURSLT[8]));
   FA1_X1_50_SVT g28772 (.A(DPATH_n_2820),
	.B(DPATH_n_2782),
	.CI(n_1301),
	.CO(n_1302),
	.S(ALURSLT[7]));
   FA1_X1_50_SVT g28773 (.A(DPATH_n_2821),
	.B(DPATH_n_2783),
	.CI(n_1300),
	.CO(n_1301),
	.S(ALURSLT[6]));
   FA1_X1_50_SVT g28774 (.A(DPATH_n_2822),
	.B(DPATH_n_2784),
	.CI(n_1299),
	.CO(n_1300),
	.S(ALURSLT[5]));
   FA1_X1_50_SVT g28775 (.A(DPATH_n_2823),
	.B(DPATH_n_2785),
	.CI(n_1298),
	.CO(n_1299),
	.S(ALURSLT[4]));
   FA1_X1_50_SVT g28776 (.A(DPATH_n_2824),
	.B(DPATH_n_2786),
	.CI(n_1297),
	.CO(n_1298),
	.S(ALURSLT[3]));
   FA1_X1_50_SVT g28777 (.A(DPATH_n_2825),
	.B(DPATH_n_2787),
	.CI(n_1296),
	.CO(n_1297),
	.S(ALURSLT[2]));
   FA1_X1_50_SVT g28778 (.A(DPATH_n_2826),
	.B(DPATH_n_2788),
	.CI(n_1295),
	.CO(n_1296),
	.S(ALURSLT[1]));
   HA1_X1_50_SVT g28779 (.A(DPATH_n_2827),
	.B(DPATH_n_2789),
	.CO(n_1295),
	.S(ALURSLT[0]));
   OAI31_X1_50_SVT g28780 (.A0(n_1153),
	.A1(n_1156),
	.A2(n_1154),
	.B0(n_1294),
	.Q(DPATH_n_2789));
   AOI222_X1_50_SVT g28781 (.A0(DPATH_n_2597),
	.A1(n_1159),
	.B0(n_1229),
	.B1(DPATH_n_2414),
	.C0(DPATH_n_2556),
	.C1(n_1251),
	.Q(n_1294));
   INV_A_OAI21_X1_50_SVT g28782 (.A0(n_1160),
	.A1N(DPATH_n_2592),
	.B0(n_1291),
	.Q(DPATH_n_2784));
   INV_A_OAI21_X1_50_SVT g28783 (.A0(n_1160),
	.A1N(DPATH_n_2593),
	.B0(n_1290),
	.Q(DPATH_n_2785));
   INV_A_OAI21_X1_50_SVT g28784 (.A0(n_1160),
	.A1N(DPATH_n_2579),
	.B0(n_1289),
	.Q(DPATH_n_2771));
   INV_A_OAI21_X1_50_SVT g28785 (.A0(n_1160),
	.A1N(DPATH_n_2568),
	.B0(n_1288),
	.Q(DPATH_n_2760));
   INV_A_OAI21_X1_50_SVT g28786 (.A0(n_1160),
	.A1N(DPATH_n_2594),
	.B0(n_1287),
	.Q(DPATH_n_2786));
   INV_A_OAI21_X1_50_SVT g28787 (.A0(n_1160),
	.A1N(DPATH_n_2595),
	.B0(n_1285),
	.Q(DPATH_n_2787));
   INV_A_OAI21_X1_50_SVT g28788 (.A0(n_1160),
	.A1N(DPATH_n_2580),
	.B0(n_1284),
	.Q(DPATH_n_2772));
   INV_A_OAI21_X1_50_SVT g28789 (.A0(n_1160),
	.A1N(DPATH_n_2596),
	.B0(n_1283),
	.Q(DPATH_n_2788));
   INV_A_OAI21_X1_50_SVT g28790 (.A0(n_1160),
	.A1N(DPATH_n_2569),
	.B0(n_1275),
	.Q(DPATH_n_2761));
   INV_A_OAI21_X1_50_SVT g28791 (.A0(n_1160),
	.A1N(DPATH_n_2581),
	.B0(n_1282),
	.Q(DPATH_n_2773));
   INV_A_OAI21_X1_50_SVT g28792 (.A0(n_1160),
	.A1N(DPATH_n_2572),
	.B0(n_1293),
	.Q(DPATH_n_2764));
   INV_A_OAI21_X1_50_SVT g28793 (.A0(n_1160),
	.A1N(DPATH_n_2573),
	.B0(n_1279),
	.Q(DPATH_n_2765));
   INV_A_OAI21_X1_50_SVT g28794 (.A0(n_1160),
	.A1N(DPATH_n_2582),
	.B0(n_1263),
	.Q(DPATH_n_2774));
   INV_A_OAI21_X1_50_SVT g28795 (.A0(n_1160),
	.A1N(DPATH_n_2574),
	.B0(n_1280),
	.Q(DPATH_n_2766));
   INV_A_OAI21_X1_50_SVT g28796 (.A0(n_1160),
	.A1N(DPATH_n_2578),
	.B0(n_1292),
	.Q(DPATH_n_2770));
   NAND2_A_NAND2_X2_50_SVT g28797 (.A0N(DPATH_n_2591),
	.A1N(n_1159),
	.B0(n_1278),
	.Q(DPATH_n_2783));
   NAND2_A_NAND2_X2_50_SVT g28798 (.A0N(DPATH_n_2584),
	.A1N(n_1159),
	.B0(n_1281),
	.Q(DPATH_n_2776));
   NAND2_A_NAND2_X2_50_SVT g28799 (.A0N(DPATH_n_2585),
	.A1N(n_1159),
	.B0(n_1276),
	.Q(DPATH_n_2777));
   NAND2_A_NAND2_X2_50_SVT g28800 (.A0N(DPATH_n_2575),
	.A1N(n_1159),
	.B0(n_1274),
	.Q(DPATH_n_2767));
   NAND2_A_NAND2_X2_50_SVT g28801 (.A0N(DPATH_n_2567),
	.A1N(n_1159),
	.B0(n_1272),
	.Q(DPATH_n_2759));
   NAND2_A_NAND2_X2_50_SVT g28802 (.A0N(DPATH_n_2586),
	.A1N(n_1159),
	.B0(n_1273),
	.Q(DPATH_n_2778));
   NAND2_A_NAND2_X2_50_SVT g28803 (.A0N(DPATH_ALU_SUM_31__624),
	.A1N(n_1159),
	.B0(n_1264),
	.Q(DPATH_n_2758));
   NAND2_A_NAND2_X2_50_SVT g28804 (.A0N(DPATH_n_2570),
	.A1N(n_1159),
	.B0(n_1271),
	.Q(DPATH_n_2762));
   NAND2_A_NAND2_X2_50_SVT g28805 (.A0N(DPATH_n_2587),
	.A1N(n_1159),
	.B0(n_1270),
	.Q(DPATH_n_2779));
   NAND2_A_NAND2_X2_50_SVT g28806 (.A0N(DPATH_n_2576),
	.A1N(n_1159),
	.B0(n_1269),
	.Q(DPATH_n_2768));
   NAND2_A_NAND2_X2_50_SVT g28807 (.A0N(DPATH_n_2588),
	.A1N(n_1159),
	.B0(n_1268),
	.Q(DPATH_n_2780));
   NAND2_A_NAND2_X2_50_SVT g28808 (.A0N(DPATH_n_2589),
	.A1N(n_1159),
	.B0(n_1267),
	.Q(DPATH_n_2781));
   NAND2_A_NAND2_X2_50_SVT g28809 (.A0N(DPATH_n_2577),
	.A1N(n_1159),
	.B0(n_1266),
	.Q(DPATH_n_2769));
   NAND2_A_NAND2_X2_50_SVT g28810 (.A0N(DPATH_n_2590),
	.A1N(n_1159),
	.B0(n_1265),
	.Q(DPATH_n_2782));
   NAND2_A_NAND2_X2_50_SVT g28811 (.A0N(DPATH_n_2571),
	.A1N(n_1159),
	.B0(n_1286),
	.Q(DPATH_n_2763));
   NAND2_A_NAND2_X2_50_SVT g28812 (.A0N(DPATH_n_2583),
	.A1N(n_1159),
	.B0(n_1277),
	.Q(DPATH_n_2775));
   AOI22_X1_50_SVT g28813 (.A0(n_1219),
	.A1(DPATH_n_2389),
	.B0(n_1247),
	.B1(DPATH_n_2506),
	.Q(n_1293));
   AOI22_X1_50_SVT g28814 (.A0(n_1227),
	.A1(DPATH_n_2395),
	.B0(n_1258),
	.B1(DPATH_n_2518),
	.Q(n_1292));
   AOI22_X1_50_SVT g28815 (.A0(n_1228),
	.A1(DPATH_n_2409),
	.B0(n_1257),
	.B1(DPATH_n_2546),
	.Q(n_1291));
   AOI22_X1_50_SVT g28816 (.A0(n_1226),
	.A1(DPATH_n_2410),
	.B0(n_1256),
	.B1(DPATH_n_2548),
	.Q(n_1290));
   AOI22_X1_50_SVT g28817 (.A0(n_1223),
	.A1(DPATH_n_2396),
	.B0(n_1246),
	.B1(DPATH_n_2520),
	.Q(n_1289));
   AOI22_X1_50_SVT g28818 (.A0(n_1218),
	.A1(DPATH_n_2385),
	.B0(n_1254),
	.B1(DPATH_n_2498),
	.Q(n_1288));
   AOI22_X1_50_SVT g28819 (.A0(n_1224),
	.A1(DPATH_n_2411),
	.B0(n_1255),
	.B1(DPATH_n_2550),
	.Q(n_1287));
   AOI22_X1_50_SVT g28820 (.A0(n_1225),
	.A1(DPATH_n_2388),
	.B0(DPATH_n_2504),
	.B1(n_1260),
	.Q(n_1286));
   AOI22_X1_50_SVT g28821 (.A0(n_1222),
	.A1(DPATH_n_2412),
	.B0(n_1245),
	.B1(DPATH_n_2552),
	.Q(n_1285));
   AOI22_X1_50_SVT g28822 (.A0(n_1220),
	.A1(DPATH_n_2397),
	.B0(n_1253),
	.B1(DPATH_n_2522),
	.Q(n_1284));
   AOI22_X1_50_SVT g28823 (.A0(n_1221),
	.A1(DPATH_n_2413),
	.B0(DPATH_n_2554),
	.B1(n_1252),
	.Q(n_1283));
   AOI22_X1_50_SVT g28824 (.A0(n_1217),
	.A1(DPATH_n_2398),
	.B0(DPATH_n_2524),
	.B1(n_1250),
	.Q(n_1282));
   AOI22_X1_50_SVT g28825 (.A0(n_1212),
	.A1(DPATH_n_2401),
	.B0(n_1244),
	.B1(DPATH_n_2530),
	.Q(n_1281));
   AOI22_X1_50_SVT g28826 (.A0(n_1211),
	.A1(DPATH_n_2391),
	.B0(n_1234),
	.B1(DPATH_n_2510),
	.Q(n_1280));
   AOI22_X1_50_SVT g28827 (.A0(n_1230),
	.A1(DPATH_n_2390),
	.B0(n_1249),
	.B1(DPATH_n_2508),
	.Q(n_1279));
   AOI22_X1_50_SVT g28828 (.A0(n_1214),
	.A1(DPATH_n_2408),
	.B0(n_1259),
	.B1(DPATH_n_2544),
	.Q(n_1278));
   AOI22_X1_50_SVT g28829 (.A0(n_1215),
	.A1(DPATH_n_2400),
	.B0(DPATH_n_2528),
	.B1(n_1243),
	.Q(n_1277));
   AOI22_X1_50_SVT g28830 (.A0(n_1209),
	.A1(DPATH_n_2402),
	.B0(DPATH_n_2532),
	.B1(n_1242),
	.Q(n_1276));
   AOI22_X1_50_SVT g28831 (.A0(n_1210),
	.A1(DPATH_n_2386),
	.B0(DPATH_n_2500),
	.B1(n_1262),
	.Q(n_1275));
   AOI22_X1_50_SVT g28832 (.A0(n_1207),
	.A1(DPATH_n_2392),
	.B0(n_1241),
	.B1(DPATH_n_2512),
	.Q(n_1274));
   AOI22_X1_50_SVT g28833 (.A0(n_1208),
	.A1(DPATH_n_2403),
	.B0(DPATH_n_2534),
	.B1(n_1240),
	.Q(n_1273));
   AOI22_X1_50_SVT g28834 (.A0(n_1199),
	.A1(DPATH_n_2384),
	.B0(n_1239),
	.B1(DPATH_n_2496),
	.Q(n_1272));
   AOI22_X1_50_SVT g28835 (.A0(n_1203),
	.A1(DPATH_n_2387),
	.B0(DPATH_n_2502),
	.B1(n_1237),
	.Q(n_1271));
   AOI22_X1_50_SVT g28836 (.A0(n_1206),
	.A1(DPATH_n_2404),
	.B0(DPATH_n_2536),
	.B1(n_1238),
	.Q(n_1270));
   AOI22_X1_50_SVT g28837 (.A0(n_1204),
	.A1(DPATH_n_2393),
	.B0(n_1236),
	.B1(DPATH_n_2514),
	.Q(n_1269));
   AOI22_X1_50_SVT g28838 (.A0(n_1205),
	.A1(DPATH_n_2405),
	.B0(DPATH_n_2538),
	.B1(n_1235),
	.Q(n_1268));
   AOI22_X1_50_SVT g28839 (.A0(n_1202),
	.A1(DPATH_n_2406),
	.B0(DPATH_n_2540),
	.B1(n_1233),
	.Q(n_1267));
   AOI22_X1_50_SVT g28840 (.A0(n_1200),
	.A1(DPATH_n_2394),
	.B0(n_1232),
	.B1(DPATH_n_2516),
	.Q(n_1266));
   AOI22_X1_50_SVT g28841 (.A0(n_1201),
	.A1(DPATH_n_2407),
	.B0(n_1231),
	.B1(DPATH_n_2542),
	.Q(n_1265));
   AOI22_X1_50_SVT g28842 (.A0(n_1216),
	.A1(DPATH_A_31_),
	.B0(n_1261),
	.B1(DPATH_B_31_),
	.Q(n_1264));
   AOI22_X1_50_SVT g28843 (.A0(n_1213),
	.A1(DPATH_n_2399),
	.B0(DPATH_n_2526),
	.B1(n_1248),
	.Q(n_1263));
   NAND2_X2_50_SVT g28844 (.A(n_1178),
	.B(n_1164),
	.Q(n_1262));
   NAND2T_X1_50_SVT g28845 (.A(n_1197),
	.B(n_1164),
	.Q(n_1261));
   NAND2T_X1_50_SVT g28846 (.A(n_1181),
	.B(n_1164),
	.Q(n_1260));
   NAND2_X2_50_SVT g28847 (.A(n_1193),
	.B(n_1164),
	.Q(n_1259));
   NAND2T_X1_50_SVT g28848 (.A(n_1196),
	.B(n_1164),
	.Q(n_1258));
   NAND2_X2_50_SVT g28849 (.A(n_1195),
	.B(n_1164),
	.Q(n_1257));
   NAND2_X2_50_SVT g28850 (.A(n_1194),
	.B(n_1164),
	.Q(n_1256));
   NAND2_X2_50_SVT g28851 (.A(n_1190),
	.B(n_1164),
	.Q(n_1255));
   NAND2_X2_50_SVT g28852 (.A(n_1182),
	.B(n_1164),
	.Q(n_1254));
   NAND2_X2_50_SVT g28853 (.A(n_1186),
	.B(n_1164),
	.Q(n_1253));
   NAND2T_X1_50_SVT g28854 (.A(n_1188),
	.B(n_1164),
	.Q(n_1252));
   NAND2T_X1_50_SVT g28855 (.A(n_1189),
	.B(n_1164),
	.Q(n_1251));
   NAND2T_X1_50_SVT g28856 (.A(n_1187),
	.B(n_1164),
	.Q(n_1250));
   NAND2_X2_50_SVT g28857 (.A(n_1180),
	.B(n_1164),
	.Q(n_1249));
   NAND2_X2_50_SVT g28858 (.A(n_1179),
	.B(n_1164),
	.Q(n_1248));
   NAND2_X2_50_SVT g28859 (.A(n_1185),
	.B(n_1164),
	.Q(n_1247));
   NAND2_X2_50_SVT g28860 (.A(n_1192),
	.B(n_1164),
	.Q(n_1246));
   NAND2T_X1_50_SVT g28861 (.A(n_1177),
	.B(n_1164),
	.Q(n_1245));
   NAND2_X2_50_SVT g28862 (.A(n_1191),
	.B(n_1164),
	.Q(n_1244));
   NAND2T_X1_50_SVT g28863 (.A(n_1184),
	.B(n_1164),
	.Q(n_1243));
   NAND2_X2_50_SVT g28864 (.A(n_1176),
	.B(n_1164),
	.Q(n_1242));
   NAND2T_X1_50_SVT g28865 (.A(n_1175),
	.B(n_1164),
	.Q(n_1241));
   NAND2_X2_50_SVT g28866 (.A(n_1174),
	.B(n_1164),
	.Q(n_1240));
   NAND2_X2_50_SVT g28867 (.A(n_1172),
	.B(n_1164),
	.Q(n_1239));
   NAND2_X2_50_SVT g28868 (.A(n_1183),
	.B(n_1164),
	.Q(n_1238));
   NAND2_X2_50_SVT g28869 (.A(n_1171),
	.B(n_1164),
	.Q(n_1237));
   NAND2T_X1_50_SVT g28870 (.A(n_1170),
	.B(n_1164),
	.Q(n_1236));
   NAND2_X2_50_SVT g28871 (.A(n_1169),
	.B(n_1164),
	.Q(n_1235));
   NAND2T_X1_50_SVT g28872 (.A(n_1167),
	.B(n_1164),
	.Q(n_1234));
   NAND2T_X1_50_SVT g28873 (.A(n_1168),
	.B(n_1164),
	.Q(n_1233));
   NAND2T_X1_50_SVT g28874 (.A(n_1173),
	.B(n_1164),
	.Q(n_1232));
   NAND2T_X1_50_SVT g28875 (.A(n_1166),
	.B(n_1164),
	.Q(n_1231));
   OAI21P2_X1_50_SVT g28876 (.A0(DPATH_n_2508),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1230));
   OAI21P2_X1_50_SVT g28877 (.A0(DPATH_n_2556),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1229));
   OAI21P2_X1_50_SVT g28878 (.A0(DPATH_n_2546),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1228));
   OAI21P2_X1_50_SVT g28879 (.A0(DPATH_n_2518),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1227));
   OAI21P2_X1_50_SVT g28880 (.A0(DPATH_n_2548),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1226));
   OAI21P2_X1_50_SVT g28881 (.A0(DPATH_n_2504),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1225));
   OAI21P2_X1_50_SVT g28882 (.A0(DPATH_n_2550),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1224));
   OAI21P2_X1_50_SVT g28883 (.A0(DPATH_n_2520),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1223));
   OAI21P2_X1_50_SVT g28884 (.A0(DPATH_n_2552),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1222));
   OAI21P2_X1_50_SVT g28885 (.A0(DPATH_n_2554),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1221));
   OAI21P2_X1_50_SVT g28886 (.A0(DPATH_n_2522),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1220));
   OAI21P2_X1_50_SVT g28887 (.A0(DPATH_n_2506),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1219));
   OAI21P2_X1_50_SVT g28888 (.A0(DPATH_n_2498),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1218));
   OAI21P2_X1_50_SVT g28889 (.A0(DPATH_n_2524),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1217));
   OAI21P2_X1_50_SVT g28890 (.A0(DPATH_B_31_),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1216));
   OAI21P2_X1_50_SVT g28891 (.A0(DPATH_n_2528),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1215));
   OAI21P2_X1_50_SVT g28892 (.A0(DPATH_n_2544),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1214));
   OAI21P2_X1_50_SVT g28893 (.A0(DPATH_n_2526),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1213));
   OAI21P2_X1_50_SVT g28894 (.A0(DPATH_n_2530),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1212));
   OAI21P2_X1_50_SVT g28895 (.A0(DPATH_n_2510),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1211));
   OAI21P2_X1_50_SVT g28896 (.A0(DPATH_n_2500),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1210));
   OAI21P2_X1_50_SVT g28897 (.A0(DPATH_n_2532),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1209));
   OAI21P2_X1_50_SVT g28898 (.A0(DPATH_n_2534),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1208));
   OAI21P2_X1_50_SVT g28899 (.A0(DPATH_n_2512),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1207));
   OAI21P2_X1_50_SVT g28900 (.A0(DPATH_n_2536),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1206));
   OAI21P2_X1_50_SVT g28901 (.A0(DPATH_n_2538),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1205));
   OAI21P2_X1_50_SVT g28902 (.A0(DPATH_n_2514),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1204));
   OAI21P2_X1_50_SVT g28903 (.A0(DPATH_n_2502),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1203));
   OAI21P2_X1_50_SVT g28904 (.A0(DPATH_n_2540),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1202));
   OAI21P2_X1_50_SVT g28905 (.A0(DPATH_n_2542),
	.A1(n_1161),
	.B0(n_1198),
	.Q(n_1201));
   OAI21P2_X1_50_SVT g28906 (.A0(DPATH_n_2516),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1200));
   OAI21P2_X1_50_SVT g28907 (.A0(DPATH_n_2496),
	.A1(n_1161),
	.B0(FE_OFN118_n_1198),
	.Q(n_1199));
   INV_A_NOR2_X2_50_SVT g28908 (.AN(DPATH_n_2532),
	.B(n_1165),
	.Q(DPATH_n_2815));
   INV_A_NOR2_X2_50_SVT g28909 (.AN(DPATH_n_2552),
	.B(n_1165),
	.Q(DPATH_n_2825));
   INV_A_NOR2_X2_50_SVT g28910 (.AN(DPATH_n_2548),
	.B(n_1165),
	.Q(DPATH_n_2823));
   INV_A_NOR2_X2_50_SVT g28911 (.AN(DPATH_n_2520),
	.B(n_1165),
	.Q(DPATH_n_2809));
   INV_A_NOR2_X2_50_SVT g28912 (.AN(DPATH_n_2550),
	.B(n_1165),
	.Q(DPATH_n_2824));
   INV_A_NOR2_X2_50_SVT g28913 (.AN(DPATH_n_2522),
	.B(n_1165),
	.Q(DPATH_n_2810));
   INV_A_NOR2_X2_50_SVT g28914 (.AN(DPATH_n_2554),
	.B(n_1165),
	.Q(DPATH_n_2826));
   INV_A_NOR2_X2_50_SVT g28915 (.AN(DPATH_n_2556),
	.B(n_1165),
	.Q(DPATH_n_2827));
   INV_A_NOR2_X2_50_SVT g28916 (.AN(DPATH_n_2524),
	.B(n_1165),
	.Q(DPATH_n_2811));
   INV_A_NOR2_X2_50_SVT g28917 (.AN(DPATH_n_2508),
	.B(n_1165),
	.Q(DPATH_n_2803));
   INV_A_NOR2_X2_50_SVT g28918 (.AN(DPATH_n_2496),
	.B(n_1165),
	.Q(DPATH_n_2797));
   INV_A_NOR2_X2_50_SVT g28919 (.AN(DPATH_n_2510),
	.B(n_1165),
	.Q(DPATH_n_2804));
   INV_A_NOR2_X2_50_SVT g28920 (.AN(DPATH_n_2506),
	.B(n_1165),
	.Q(DPATH_n_2802));
   INV_A_NOR2_X2_50_SVT g28921 (.AN(DPATH_n_2528),
	.B(n_1165),
	.Q(DPATH_n_2813));
   INV_A_NOR2_X2_50_SVT g28922 (.AN(DPATH_n_2500),
	.B(n_1165),
	.Q(DPATH_n_2799));
   INV_A_NOR2_X2_50_SVT g28923 (.AN(DPATH_n_2526),
	.B(n_1165),
	.Q(DPATH_n_2812));
   INV_A_NOR2_X2_50_SVT g28924 (.AN(DPATH_n_2518),
	.B(n_1165),
	.Q(DPATH_n_2808));
   INV_A_NOR2_X2_50_SVT g28925 (.AN(DPATH_n_2512),
	.B(n_1165),
	.Q(DPATH_n_2805));
   INV_A_NOR2_X2_50_SVT g28926 (.AN(DPATH_n_2534),
	.B(n_1165),
	.Q(DPATH_n_2816));
   INV_A_NOR2_X2_50_SVT g28927 (.AN(DPATH_n_2498),
	.B(n_1165),
	.Q(DPATH_n_2798));
   INV_A_NOR2_X2_50_SVT g28928 (.AN(DPATH_n_2502),
	.B(n_1165),
	.Q(DPATH_n_2800));
   INV_A_NOR2_X2_50_SVT g28929 (.AN(DPATH_n_2536),
	.B(n_1165),
	.Q(DPATH_n_2817));
   INV_A_NOR2_X2_50_SVT g28930 (.AN(DPATH_n_2514),
	.B(n_1165),
	.Q(DPATH_n_2806));
   INV_A_NOR2_X2_50_SVT g28931 (.AN(DPATH_n_2538),
	.B(n_1165),
	.Q(DPATH_n_2818));
   INV_A_NOR2_X2_50_SVT g28932 (.AN(DPATH_n_2540),
	.B(n_1165),
	.Q(DPATH_n_2819));
   INV_A_NOR2_X2_50_SVT g28933 (.AN(DPATH_n_2530),
	.B(n_1165),
	.Q(DPATH_n_2814));
   INV_A_NOR2_X2_50_SVT g28934 (.AN(DPATH_B_31_),
	.B(n_1165),
	.Q(DPATH_n_2796));
   INV_A_NOR2_X2_50_SVT g28935 (.AN(DPATH_n_2516),
	.B(n_1165),
	.Q(DPATH_n_2807));
   INV_A_NOR2_X2_50_SVT g28936 (.AN(DPATH_n_2542),
	.B(n_1165),
	.Q(DPATH_n_2820));
   INV_A_NOR2_X2_50_SVT g28937 (.AN(DPATH_n_2546),
	.B(n_1165),
	.Q(DPATH_n_2822));
   INV_A_NOR2_X2_50_SVT g28938 (.AN(DPATH_n_2504),
	.B(n_1165),
	.Q(DPATH_n_2801));
   INV_A_NOR2_X2_50_SVT g28939 (.AN(DPATH_n_2544),
	.B(n_1165),
	.Q(DPATH_n_2821));
   MUXI2_X1_50_SVT g28940 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1197),
	.S0(DPATH_A_31_));
   MUXI2_X1_50_SVT g28941 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1196),
	.S0(DPATH_n_2395));
   MUXI2_X1_50_SVT g28942 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1195),
	.S0(DPATH_n_2409));
   MUXI2_X1_50_SVT g28943 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1194),
	.S0(DPATH_n_2410));
   MUXI2_X1_50_SVT g28944 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1193),
	.S0(DPATH_n_2408));
   MUXI2_X1_50_SVT g28945 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1192),
	.S0(DPATH_n_2396));
   MUXI2_X1_50_SVT g28946 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1191),
	.S0(DPATH_n_2401));
   MUXI2_X1_50_SVT g28947 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1190),
	.S0(DPATH_n_2411));
   MUXI2_X1_50_SVT g28948 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1189),
	.S0(DPATH_n_2414));
   MUXI2_X1_50_SVT g28949 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1188),
	.S0(DPATH_n_2413));
   MUXI2_X1_50_SVT g28950 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1187),
	.S0(DPATH_n_2398));
   MUXI2_X1_50_SVT g28951 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1186),
	.S0(DPATH_n_2397));
   MUXI2_X1_50_SVT g28952 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1185),
	.S0(DPATH_n_2389));
   MUXI2_X1_50_SVT g28953 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1184),
	.S0(DPATH_n_2400));
   MUXI2_X1_50_SVT g28954 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1183),
	.S0(DPATH_n_2404));
   MUXI2_X1_50_SVT g28955 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1182),
	.S0(DPATH_n_2385));
   MUXI2_X1_50_SVT g28956 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1181),
	.S0(DPATH_n_2388));
   MUXI2_X1_50_SVT g28957 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1180),
	.S0(DPATH_n_2390));
   MUXI2_X1_50_SVT g28958 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1179),
	.S0(DPATH_n_2399));
   MUXI2_X1_50_SVT g28959 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1178),
	.S0(DPATH_n_2386));
   MUXI2_X1_50_SVT g28960 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1177),
	.S0(DPATH_n_2412));
   MUXI2_X1_50_SVT g28961 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1176),
	.S0(DPATH_n_2402));
   MUXI2_X1_50_SVT g28962 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1175),
	.S0(DPATH_n_2392));
   MUXI2_X1_50_SVT g28963 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1174),
	.S0(DPATH_n_2403));
   MUXI2_X1_50_SVT g28964 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1173),
	.S0(DPATH_n_2394));
   MUXI2_X1_50_SVT g28965 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1172),
	.S0(DPATH_n_2384));
   MUXI2_X1_50_SVT g28966 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1171),
	.S0(DPATH_n_2387));
   MUXI2_X1_50_SVT g28967 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1170),
	.S0(DPATH_n_2393));
   MUXI2_X1_50_SVT g28968 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1169),
	.S0(DPATH_n_2405));
   MUXI2_X1_50_SVT g28969 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1168),
	.S0(DPATH_n_2406));
   MUXI2_X1_50_SVT g28970 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1167),
	.S0(DPATH_n_2391));
   MUXI2_X1_50_SVT g28971 (.A(FE_OFN24_n_1162),
	.B(n_1158),
	.Q(n_1166),
	.S0(DPATH_n_2407));
   NOR2P3_X2_50_SVT g28972 (.A(n_1163),
	.B(n_1148),
	.Q(n_1198));
   CLKINV_X4_50_SVT g28975 (.A(n_1163),
	.Q(n_1164));
   INV_A_NOR2_X0_50_SVT g28977 (.AN(n_1155),
	.B(n_1156),
	.Q(n_1163));
   NOR2_X0_50_SVT g28978 (.A(n_1154),
	.B(n_1157),
	.Q(n_1162));
   INV_X2_50_SVT g28979 (.A(n_1160),
	.Q(n_1159));
   CLKNAND2_X2_50_SVT g28981 (.A(n_1157),
	.B(n_1147),
	.Q(n_1160));
   CLKAND2_X2_50_SVT g28982 (.A(n_1156),
	.B(n_1154),
	.Q(n_1158));
   OAI221_X0_50_SVT g28984 (.A0(INSTR[12]),
	.A1(n_1147),
	.B0(INSTR[4]),
	.B1(n_2706),
	.C0(n_1152),
	.Q(n_1157));
   INV_A_NOR2_X0_50_SVT g28985 (.AN(INSTR[14]),
	.B(n_1147),
	.Q(n_1155));
   OR2_X1_50_SVT g28986 (.A(n_1147),
	.B(INSTR[14]),
	.Q(n_1154));
   AOI22_X1_50_SVT g28988 (.A0(n_1150),
	.A1(DPATH_A_31_),
	.B0(DPATH_ALU_SUM_31__624),
	.B1(n_1149),
	.Q(n_1153));
   INV_A_NAND3_X0_50_SVT g28989 (.AN(n_2708),
	.B(INSTR[30]),
	.C(n_1151),
	.Q(n_1152));
   NOR3_X0_50_SVT g28991 (.A(INSTR[14]),
	.B(INSTR[13]),
	.C(INSTR[12]),
	.Q(n_1151));
   INV_A_NAND2_X2_50_SVT g28992 (.AN(DPATH_ALU_SUM_31__624),
	.B(DPATH_B_31_),
	.Q(n_1150));
   INV_A_NOR2_X0_50_SVT g79924 (.AN(n_1158),
	.B(n_1155),
	.Q(n_1148));
   INV_A_NAND2_X2_50_SVT g28995 (.AN(n_1151),
	.B(INSTR[4]),
	.Q(n_1147));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_0_ (.CK(CTS_5),
	.D(PC[0]),
	.Q(PC[0]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_1_ (.CK(CTS_6),
	.D(n_40),
	.Q(PC[1]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_2_ (.CK(CTS_5),
	.D(n_44),
	.Q(PC[2]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_3_ (.CK(CTS_5),
	.D(n_41),
	.Q(PC[3]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_4_ (.CK(CTS_5),
	.D(n_42),
	.Q(PC[4]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_5_ (.CK(CTS_5),
	.D(n_32),
	.Q(PC[5]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_6_ (.CK(CTS_5),
	.D(n_51),
	.Q(PC[6]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_7_ (.CK(CTS_5),
	.D(n_50),
	.Q(PC[7]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_8_ (.CK(CTS_5),
	.D(n_45),
	.Q(PC[8]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_9_ (.CK(CTS_6),
	.D(n_48),
	.Q(PC[9]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_10_ (.CK(CTS_6),
	.D(n_49),
	.Q(PC[10]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_11_ (.CK(CTS_6),
	.D(n_60),
	.Q(PC[11]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_12_ (.CK(CTS_6),
	.D(n_52),
	.Q(PC[12]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_13_ (.CK(CTS_6),
	.D(n_56),
	.Q(PC[13]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_14_ (.CK(CTS_6),
	.D(n_38),
	.Q(PC[14]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_15_ (.CK(CTS_6),
	.D(n_35),
	.Q(PC[15]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_16_ (.CK(CTS_6),
	.D(n_43),
	.Q(PC[16]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_17_ (.CK(CTS_9),
	.D(n_47),
	.Q(PC[17]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_18_ (.CK(CTS_6),
	.D(n_29),
	.Q(PC[18]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_19_ (.CK(CTS_6),
	.D(n_36),
	.Q(PC[19]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_20_ (.CK(CTS_6),
	.D(n_31),
	.Q(PC[20]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_21_ (.CK(CTS_6),
	.D(n_39),
	.Q(PC[21]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_22_ (.CK(CTS_6),
	.D(n_57),
	.Q(PC[22]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_23_ (.CK(CTS_6),
	.D(n_55),
	.Q(PC[23]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_24_ (.CK(CTS_6),
	.D(n_33),
	.Q(PC[24]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_25_ (.CK(CTS_6),
	.D(n_54),
	.Q(PC[25]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_26_ (.CK(CTS_6),
	.D(n_46),
	.Q(PC[26]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_27_ (.CK(CTS_2),
	.D(n_34),
	.Q(PC[27]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_28_ (.CK(CTS_2),
	.D(n_30),
	.Q(PC[28]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_29_ (.CK(CTS_2),
	.D(n_37),
	.Q(PC[29]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_30_ (.CK(CTS_2),
	.D(n_59),
	.Q(PC[30]),
	.RN(n_2672));
   DFFRQ_X2_50_SVT DPATH_PCREG_Q_reg_31_ (.CK(CTS_2),
	.D(n_58),
	.Q(PC[31]),
	.RN(n_2672));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__0_ (.CK(CTS_15),
	.D(n_389),
	.Q(DPATH_RF_MEMORY_1__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__1_ (.CK(CTS_16),
	.D(n_374),
	.Q(DPATH_RF_MEMORY_1__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__2_ (.CK(CTS_11),
	.D(n_161),
	.Q(DPATH_RF_MEMORY_1__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__3_ (.CK(CTS_61),
	.D(n_402),
	.Q(DPATH_RF_MEMORY_1__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__4_ (.CK(CTS_10),
	.D(n_372),
	.Q(DPATH_RF_MEMORY_1__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__5_ (.CK(CTS_11),
	.D(n_371),
	.Q(DPATH_RF_MEMORY_1__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__6_ (.CK(CTS_50),
	.D(n_369),
	.Q(DPATH_RF_MEMORY_1__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__7_ (.CK(CTS_19),
	.D(n_368),
	.Q(DPATH_RF_MEMORY_1__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__8_ (.CK(CTS_61),
	.D(n_367),
	.Q(DPATH_RF_MEMORY_1__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__9_ (.CK(CTS_23),
	.D(n_364),
	.Q(DPATH_RF_MEMORY_1__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__10_ (.CK(CTS_14),
	.D(n_354),
	.Q(DPATH_RF_MEMORY_1__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__11_ (.CK(CTS_54),
	.D(n_356),
	.Q(DPATH_RF_MEMORY_1__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__12_ (.CK(CTS_44),
	.D(n_335),
	.Q(DPATH_RF_MEMORY_1__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__13_ (.CK(CTS_11),
	.D(n_350),
	.Q(DPATH_RF_MEMORY_1__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__14_ (.CK(CTS_47),
	.D(n_340),
	.Q(DPATH_RF_MEMORY_1__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__15_ (.CK(CTS_37),
	.D(n_333),
	.Q(DPATH_RF_MEMORY_1__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__16_ (.CK(CTS_56),
	.D(n_328),
	.Q(DPATH_RF_MEMORY_1__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__17_ (.CK(CTS_57),
	.D(n_327),
	.Q(DPATH_RF_MEMORY_1__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__18_ (.CK(CTS_37),
	.D(n_326),
	.Q(DPATH_RF_MEMORY_1__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__19_ (.CK(CTS_37),
	.D(n_325),
	.Q(DPATH_RF_MEMORY_1__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__20_ (.CK(CTS_30),
	.D(n_324),
	.Q(DPATH_RF_MEMORY_1__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__21_ (.CK(CTS_56),
	.D(n_323),
	.Q(DPATH_RF_MEMORY_1__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__22_ (.CK(CTS_56),
	.D(n_322),
	.Q(DPATH_RF_MEMORY_1__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__23_ (.CK(CTS_34),
	.D(n_321),
	.Q(DPATH_RF_MEMORY_1__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__24_ (.CK(CTS_56),
	.D(n_320),
	.Q(DPATH_RF_MEMORY_1__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__25_ (.CK(CTS_57),
	.D(n_319),
	.Q(DPATH_RF_MEMORY_1__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__26_ (.CK(CTS_44),
	.D(n_315),
	.Q(DPATH_RF_MEMORY_1__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__27_ (.CK(CTS_36),
	.D(n_318),
	.Q(DPATH_RF_MEMORY_1__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__28_ (.CK(CTS_29),
	.D(n_317),
	.Q(DPATH_RF_MEMORY_1__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__29_ (.CK(CTS_56),
	.D(n_316),
	.Q(DPATH_RF_MEMORY_1__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__30_ (.CK(CTS_56),
	.D(n_314),
	.Q(DPATH_RF_MEMORY_1__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_1__31_ (.CK(CTS_36),
	.D(n_313),
	.Q(DPATH_RF_MEMORY_1__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__0_ (.CK(CTS_15),
	.D(n_588),
	.Q(DPATH_RF_MEMORY_2__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__1_ (.CK(CTS_16),
	.D(n_587),
	.Q(DPATH_RF_MEMORY_2__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__2_ (.CK(CTS_11),
	.D(n_167),
	.Q(DPATH_RF_MEMORY_2__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__3_ (.CK(CTS_61),
	.D(n_585),
	.Q(DPATH_RF_MEMORY_2__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__4_ (.CK(CTS_10),
	.D(n_586),
	.Q(DPATH_RF_MEMORY_2__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__5_ (.CK(CTS_11),
	.D(n_584),
	.Q(DPATH_RF_MEMORY_2__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__6_ (.CK(CTS_50),
	.D(n_583),
	.Q(DPATH_RF_MEMORY_2__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__7_ (.CK(CTS_19),
	.D(n_582),
	.Q(DPATH_RF_MEMORY_2__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__8_ (.CK(CTS_61),
	.D(n_581),
	.Q(DPATH_RF_MEMORY_2__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__9_ (.CK(CTS_61),
	.D(n_580),
	.Q(DPATH_RF_MEMORY_2__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__10_ (.CK(CTS_14),
	.D(n_579),
	.Q(DPATH_RF_MEMORY_2__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__11_ (.CK(CTS_54),
	.D(n_578),
	.Q(DPATH_RF_MEMORY_2__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__12_ (.CK(CTS_44),
	.D(n_577),
	.Q(DPATH_RF_MEMORY_2__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__13_ (.CK(CTS_11),
	.D(n_576),
	.Q(DPATH_RF_MEMORY_2__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__14_ (.CK(CTS_53),
	.D(n_575),
	.Q(DPATH_RF_MEMORY_2__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__15_ (.CK(CTS_37),
	.D(n_574),
	.Q(DPATH_RF_MEMORY_2__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__16_ (.CK(CTS_56),
	.D(n_573),
	.Q(DPATH_RF_MEMORY_2__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__17_ (.CK(CTS_57),
	.D(n_572),
	.Q(DPATH_RF_MEMORY_2__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__18_ (.CK(CTS_37),
	.D(n_570),
	.Q(DPATH_RF_MEMORY_2__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__19_ (.CK(CTS_37),
	.D(n_569),
	.Q(DPATH_RF_MEMORY_2__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__20_ (.CK(CTS_30),
	.D(n_571),
	.Q(DPATH_RF_MEMORY_2__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__21_ (.CK(CTS_56),
	.D(n_568),
	.Q(DPATH_RF_MEMORY_2__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__22_ (.CK(CTS_56),
	.D(n_567),
	.Q(DPATH_RF_MEMORY_2__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__23_ (.CK(CTS_36),
	.D(n_566),
	.Q(DPATH_RF_MEMORY_2__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__24_ (.CK(CTS_56),
	.D(n_565),
	.Q(DPATH_RF_MEMORY_2__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__25_ (.CK(CTS_57),
	.D(n_564),
	.Q(DPATH_RF_MEMORY_2__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__26_ (.CK(CTS_44),
	.D(n_563),
	.Q(DPATH_RF_MEMORY_2__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__27_ (.CK(CTS_36),
	.D(n_562),
	.Q(DPATH_RF_MEMORY_2__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__28_ (.CK(CTS_17),
	.D(n_561),
	.Q(DPATH_RF_MEMORY_2__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__29_ (.CK(CTS_56),
	.D(n_560),
	.Q(DPATH_RF_MEMORY_2__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__30_ (.CK(CTS_56),
	.D(n_559),
	.Q(DPATH_RF_MEMORY_2__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_2__31_ (.CK(CTS_36),
	.D(n_558),
	.Q(DPATH_RF_MEMORY_2__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__0_ (.CK(CTS_15),
	.D(n_280),
	.Q(DPATH_RF_MEMORY_3__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__1_ (.CK(CTS_50),
	.D(n_279),
	.Q(DPATH_RF_MEMORY_3__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__2_ (.CK(CTS_11),
	.D(n_158),
	.Q(DPATH_RF_MEMORY_3__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__3_ (.CK(CTS_19),
	.D(n_277),
	.Q(DPATH_RF_MEMORY_3__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__4_ (.CK(CTS_10),
	.D(n_278),
	.Q(DPATH_RF_MEMORY_3__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__5_ (.CK(CTS_40),
	.D(n_276),
	.Q(DPATH_RF_MEMORY_3__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__6_ (.CK(CTS_16),
	.D(n_275),
	.Q(DPATH_RF_MEMORY_3__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__7_ (.CK(CTS_19),
	.D(n_274),
	.Q(DPATH_RF_MEMORY_3__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__8_ (.CK(CTS_19),
	.D(n_273),
	.Q(DPATH_RF_MEMORY_3__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__9_ (.CK(CTS_19),
	.D(n_272),
	.Q(DPATH_RF_MEMORY_3__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__10_ (.CK(CTS_41),
	.D(n_271),
	.Q(DPATH_RF_MEMORY_3__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__11_ (.CK(CTS_28),
	.D(n_270),
	.Q(DPATH_RF_MEMORY_3__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__12_ (.CK(CTS_59),
	.D(n_268),
	.Q(DPATH_RF_MEMORY_3__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__13_ (.CK(CTS_14),
	.D(n_266),
	.Q(DPATH_RF_MEMORY_3__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__14_ (.CK(CTS_53),
	.D(n_262),
	.Q(DPATH_RF_MEMORY_3__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__15_ (.CK(CTS_37),
	.D(n_260),
	.Q(DPATH_RF_MEMORY_3__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__16_ (.CK(CTS_53),
	.D(n_257),
	.Q(DPATH_RF_MEMORY_3__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__17_ (.CK(CTS_38),
	.D(n_253),
	.Q(DPATH_RF_MEMORY_3__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__18_ (.CK(CTS_37),
	.D(n_251),
	.Q(DPATH_RF_MEMORY_3__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__19_ (.CK(CTS_37),
	.D(n_244),
	.Q(DPATH_RF_MEMORY_3__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__20_ (.CK(CTS_30),
	.D(n_242),
	.Q(DPATH_RF_MEMORY_3__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__21_ (.CK(CTS_53),
	.D(n_240),
	.Q(DPATH_RF_MEMORY_3__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__22_ (.CK(CTS_53),
	.D(n_236),
	.Q(DPATH_RF_MEMORY_3__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__23_ (.CK(CTS_36),
	.D(n_234),
	.Q(DPATH_RF_MEMORY_3__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__24_ (.CK(CTS_55),
	.D(n_232),
	.Q(DPATH_RF_MEMORY_3__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__25_ (.CK(CTS_57),
	.D(n_228),
	.Q(DPATH_RF_MEMORY_3__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__26_ (.CK(CTS_59),
	.D(n_225),
	.Q(DPATH_RF_MEMORY_3__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__27_ (.CK(CTS_35),
	.D(n_223),
	.Q(DPATH_RF_MEMORY_3__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__28_ (.CK(CTS_29),
	.D(n_220),
	.Q(DPATH_RF_MEMORY_3__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__29_ (.CK(CTS_55),
	.D(n_219),
	.Q(DPATH_RF_MEMORY_3__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__30_ (.CK(CTS_53),
	.D(n_218),
	.Q(DPATH_RF_MEMORY_3__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_3__31_ (.CK(CTS_36),
	.D(n_217),
	.Q(DPATH_RF_MEMORY_3__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__0_ (.CK(CTS_19),
	.D(n_769),
	.Q(DPATH_RF_MEMORY_4__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__1_ (.CK(CTS_50),
	.D(n_757),
	.Q(DPATH_RF_MEMORY_4__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__2_ (.CK(CTS_11),
	.D(n_172),
	.Q(DPATH_RF_MEMORY_4__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__3_ (.CK(CTS_22),
	.D(n_760),
	.Q(DPATH_RF_MEMORY_4__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__4_ (.CK(CTS_36),
	.D(n_756),
	.Q(DPATH_RF_MEMORY_4__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__5_ (.CK(CTS_40),
	.D(n_751),
	.Q(DPATH_RF_MEMORY_4__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__6_ (.CK(CTS_16),
	.D(n_750),
	.Q(DPATH_RF_MEMORY_4__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__7_ (.CK(CTS_19),
	.D(n_747),
	.Q(DPATH_RF_MEMORY_4__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__8_ (.CK(CTS_19),
	.D(n_744),
	.Q(DPATH_RF_MEMORY_4__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__9_ (.CK(CTS_19),
	.D(n_740),
	.Q(DPATH_RF_MEMORY_4__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__10_ (.CK(CTS_14),
	.D(n_738),
	.Q(DPATH_RF_MEMORY_4__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__11_ (.CK(CTS_28),
	.D(n_735),
	.Q(DPATH_RF_MEMORY_4__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__12_ (.CK(CTS_30),
	.D(n_734),
	.Q(DPATH_RF_MEMORY_4__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__13_ (.CK(CTS_14),
	.D(n_733),
	.Q(DPATH_RF_MEMORY_4__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__14_ (.CK(CTS_45),
	.D(n_732),
	.Q(DPATH_RF_MEMORY_4__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__15_ (.CK(CTS_37),
	.D(n_731),
	.Q(DPATH_RF_MEMORY_4__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__16_ (.CK(CTS_45),
	.D(n_730),
	.Q(DPATH_RF_MEMORY_4__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__17_ (.CK(CTS_38),
	.D(n_728),
	.Q(DPATH_RF_MEMORY_4__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__18_ (.CK(CTS_37),
	.D(n_727),
	.Q(DPATH_RF_MEMORY_4__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__19_ (.CK(CTS_37),
	.D(n_729),
	.Q(DPATH_RF_MEMORY_4__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__20_ (.CK(CTS_30),
	.D(n_726),
	.Q(DPATH_RF_MEMORY_4__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__21_ (.CK(CTS_52),
	.D(n_725),
	.Q(DPATH_RF_MEMORY_4__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__22_ (.CK(CTS_53),
	.D(n_724),
	.Q(DPATH_RF_MEMORY_4__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__23_ (.CK(CTS_36),
	.D(n_722),
	.Q(DPATH_RF_MEMORY_4__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__24_ (.CK(CTS_55),
	.D(n_721),
	.Q(DPATH_RF_MEMORY_4__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__25_ (.CK(CTS_38),
	.D(n_720),
	.Q(DPATH_RF_MEMORY_4__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__26_ (.CK(CTS_43),
	.D(n_719),
	.Q(DPATH_RF_MEMORY_4__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__27_ (.CK(CTS_36),
	.D(n_718),
	.Q(DPATH_RF_MEMORY_4__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__28_ (.CK(CTS_59),
	.D(n_715),
	.Q(DPATH_RF_MEMORY_4__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__29_ (.CK(CTS_52),
	.D(n_712),
	.Q(DPATH_RF_MEMORY_4__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__30_ (.CK(CTS_53),
	.D(n_710),
	.Q(DPATH_RF_MEMORY_4__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_4__31_ (.CK(CTS_36),
	.D(n_708),
	.Q(DPATH_RF_MEMORY_4__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__0_ (.CK(CTS_61),
	.D(n_490),
	.Q(DPATH_RF_MEMORY_5__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__1_ (.CK(CTS_50),
	.D(n_488),
	.Q(DPATH_RF_MEMORY_5__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__2_ (.CK(CTS_14),
	.D(n_165),
	.Q(DPATH_RF_MEMORY_5__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__3_ (.CK(CTS_61),
	.D(n_489),
	.Q(DPATH_RF_MEMORY_5__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__4_ (.CK(CTS_32),
	.D(n_487),
	.Q(DPATH_RF_MEMORY_5__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__5_ (.CK(CTS_40),
	.D(n_486),
	.Q(DPATH_RF_MEMORY_5__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__6_ (.CK(CTS_50),
	.D(n_485),
	.Q(DPATH_RF_MEMORY_5__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__7_ (.CK(CTS_61),
	.D(n_484),
	.Q(DPATH_RF_MEMORY_5__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__8_ (.CK(CTS_61),
	.D(n_483),
	.Q(DPATH_RF_MEMORY_5__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__9_ (.CK(CTS_23),
	.D(n_482),
	.Q(DPATH_RF_MEMORY_5__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__10_ (.CK(CTS_40),
	.D(n_481),
	.Q(DPATH_RF_MEMORY_5__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__11_ (.CK(CTS_55),
	.D(n_480),
	.Q(DPATH_RF_MEMORY_5__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__12_ (.CK(CTS_44),
	.D(n_477),
	.Q(DPATH_RF_MEMORY_5__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__13_ (.CK(CTS_14),
	.D(n_474),
	.Q(DPATH_RF_MEMORY_5__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__14_ (.CK(CTS_53),
	.D(n_472),
	.Q(DPATH_RF_MEMORY_5__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__15_ (.CK(CTS_37),
	.D(n_470),
	.Q(DPATH_RF_MEMORY_5__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__16_ (.CK(CTS_53),
	.D(n_466),
	.Q(DPATH_RF_MEMORY_5__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__17_ (.CK(CTS_57),
	.D(n_545),
	.Q(DPATH_RF_MEMORY_5__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__18_ (.CK(CTS_37),
	.D(n_557),
	.Q(DPATH_RF_MEMORY_5__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__19_ (.CK(CTS_37),
	.D(n_551),
	.Q(DPATH_RF_MEMORY_5__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__20_ (.CK(CTS_30),
	.D(n_549),
	.Q(DPATH_RF_MEMORY_5__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__21_ (.CK(CTS_56),
	.D(n_543),
	.Q(DPATH_RF_MEMORY_5__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__22_ (.CK(CTS_56),
	.D(n_541),
	.Q(DPATH_RF_MEMORY_5__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__23_ (.CK(CTS_36),
	.D(n_539),
	.Q(DPATH_RF_MEMORY_5__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__24_ (.CK(CTS_56),
	.D(n_535),
	.Q(DPATH_RF_MEMORY_5__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__25_ (.CK(CTS_57),
	.D(n_532),
	.Q(DPATH_RF_MEMORY_5__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__26_ (.CK(CTS_44),
	.D(n_530),
	.Q(DPATH_RF_MEMORY_5__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__27_ (.CK(CTS_36),
	.D(n_527),
	.Q(DPATH_RF_MEMORY_5__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__28_ (.CK(CTS_4),
	.D(n_525),
	.Q(DPATH_RF_MEMORY_5__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__29_ (.CK(CTS_55),
	.D(n_524),
	.Q(DPATH_RF_MEMORY_5__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__30_ (.CK(CTS_56),
	.D(n_523),
	.Q(DPATH_RF_MEMORY_5__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_5__31_ (.CK(CTS_32),
	.D(n_522),
	.Q(DPATH_RF_MEMORY_5__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__0_ (.CK(CTS_61),
	.D(n_681),
	.Q(DPATH_RF_MEMORY_6__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__1_ (.CK(CTS_50),
	.D(n_680),
	.Q(DPATH_RF_MEMORY_6__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__2_ (.CK(CTS_11),
	.D(n_170),
	.Q(DPATH_RF_MEMORY_6__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__3_ (.CK(CTS_61),
	.D(n_679),
	.Q(DPATH_RF_MEMORY_6__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__4_ (.CK(CTS_36),
	.D(n_678),
	.Q(DPATH_RF_MEMORY_6__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__5_ (.CK(CTS_40),
	.D(n_677),
	.Q(DPATH_RF_MEMORY_6__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__6_ (.CK(CTS_61),
	.D(n_676),
	.Q(DPATH_RF_MEMORY_6__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__7_ (.CK(CTS_61),
	.D(n_675),
	.Q(DPATH_RF_MEMORY_6__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__8_ (.CK(CTS_61),
	.D(n_674),
	.Q(DPATH_RF_MEMORY_6__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__9_ (.CK(CTS_61),
	.D(n_673),
	.Q(DPATH_RF_MEMORY_6__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__10_ (.CK(CTS_11),
	.D(n_672),
	.Q(DPATH_RF_MEMORY_6__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__11_ (.CK(CTS_55),
	.D(n_671),
	.Q(DPATH_RF_MEMORY_6__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__12_ (.CK(CTS_44),
	.D(n_670),
	.Q(DPATH_RF_MEMORY_6__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__13_ (.CK(CTS_11),
	.D(n_669),
	.Q(DPATH_RF_MEMORY_6__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__14_ (.CK(CTS_53),
	.D(n_668),
	.Q(DPATH_RF_MEMORY_6__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__15_ (.CK(CTS_37),
	.D(n_667),
	.Q(DPATH_RF_MEMORY_6__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__16_ (.CK(CTS_53),
	.D(n_665),
	.Q(DPATH_RF_MEMORY_6__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__17_ (.CK(CTS_38),
	.D(n_664),
	.Q(DPATH_RF_MEMORY_6__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__18_ (.CK(CTS_37),
	.D(n_666),
	.Q(DPATH_RF_MEMORY_6__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__19_ (.CK(CTS_38),
	.D(n_663),
	.Q(DPATH_RF_MEMORY_6__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__20_ (.CK(CTS_30),
	.D(n_662),
	.Q(DPATH_RF_MEMORY_6__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__21_ (.CK(CTS_53),
	.D(n_661),
	.Q(DPATH_RF_MEMORY_6__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__22_ (.CK(CTS_56),
	.D(n_660),
	.Q(DPATH_RF_MEMORY_6__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__23_ (.CK(CTS_32),
	.D(n_659),
	.Q(DPATH_RF_MEMORY_6__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__24_ (.CK(CTS_55),
	.D(n_658),
	.Q(DPATH_RF_MEMORY_6__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__25_ (.CK(CTS_57),
	.D(n_657),
	.Q(DPATH_RF_MEMORY_6__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__26_ (.CK(CTS_44),
	.D(n_656),
	.Q(DPATH_RF_MEMORY_6__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__27_ (.CK(CTS_36),
	.D(n_655),
	.Q(DPATH_RF_MEMORY_6__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__28_ (.CK(CTS_4),
	.D(n_654),
	.Q(DPATH_RF_MEMORY_6__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__29_ (.CK(CTS_55),
	.D(n_653),
	.Q(DPATH_RF_MEMORY_6__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__30_ (.CK(CTS_56),
	.D(n_652),
	.Q(DPATH_RF_MEMORY_6__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_6__31_ (.CK(CTS_36),
	.D(n_651),
	.Q(DPATH_RF_MEMORY_6__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__0_ (.CK(CTS_19),
	.D(n_433),
	.Q(DPATH_RF_MEMORY_7__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__1_ (.CK(CTS_50),
	.D(n_431),
	.Q(DPATH_RF_MEMORY_7__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__2_ (.CK(CTS_11),
	.D(n_162),
	.Q(DPATH_RF_MEMORY_7__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__3_ (.CK(CTS_61),
	.D(n_432),
	.Q(DPATH_RF_MEMORY_7__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__4_ (.CK(CTS_32),
	.D(n_429),
	.Q(DPATH_RF_MEMORY_7__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__5_ (.CK(CTS_11),
	.D(n_430),
	.Q(DPATH_RF_MEMORY_7__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__6_ (.CK(CTS_50),
	.D(n_428),
	.Q(DPATH_RF_MEMORY_7__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__7_ (.CK(CTS_19),
	.D(n_427),
	.Q(DPATH_RF_MEMORY_7__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__8_ (.CK(CTS_19),
	.D(n_426),
	.Q(DPATH_RF_MEMORY_7__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__9_ (.CK(CTS_19),
	.D(n_425),
	.Q(DPATH_RF_MEMORY_7__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__10_ (.CK(CTS_40),
	.D(n_424),
	.Q(DPATH_RF_MEMORY_7__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__11_ (.CK(CTS_52),
	.D(n_423),
	.Q(DPATH_RF_MEMORY_7__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__12_ (.CK(CTS_44),
	.D(n_421),
	.Q(DPATH_RF_MEMORY_7__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__13_ (.CK(CTS_11),
	.D(n_422),
	.Q(DPATH_RF_MEMORY_7__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__14_ (.CK(CTS_53),
	.D(n_420),
	.Q(DPATH_RF_MEMORY_7__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__15_ (.CK(CTS_38),
	.D(n_419),
	.Q(DPATH_RF_MEMORY_7__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__16_ (.CK(CTS_53),
	.D(n_418),
	.Q(DPATH_RF_MEMORY_7__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__17_ (.CK(CTS_57),
	.D(n_417),
	.Q(DPATH_RF_MEMORY_7__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__18_ (.CK(CTS_38),
	.D(n_415),
	.Q(DPATH_RF_MEMORY_7__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__19_ (.CK(CTS_38),
	.D(n_416),
	.Q(DPATH_RF_MEMORY_7__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__20_ (.CK(CTS_30),
	.D(n_413),
	.Q(DPATH_RF_MEMORY_7__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__21_ (.CK(CTS_53),
	.D(n_414),
	.Q(DPATH_RF_MEMORY_7__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__22_ (.CK(CTS_56),
	.D(n_412),
	.Q(DPATH_RF_MEMORY_7__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__23_ (.CK(CTS_32),
	.D(n_411),
	.Q(DPATH_RF_MEMORY_7__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__24_ (.CK(CTS_56),
	.D(n_410),
	.Q(DPATH_RF_MEMORY_7__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__25_ (.CK(CTS_57),
	.D(n_409),
	.Q(DPATH_RF_MEMORY_7__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__26_ (.CK(CTS_44),
	.D(n_408),
	.Q(DPATH_RF_MEMORY_7__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__27_ (.CK(CTS_8),
	.D(n_407),
	.Q(DPATH_RF_MEMORY_7__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__28_ (.CK(CTS_17),
	.D(n_406),
	.Q(DPATH_RF_MEMORY_7__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__29_ (.CK(CTS_55),
	.D(n_405),
	.Q(DPATH_RF_MEMORY_7__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__30_ (.CK(CTS_56),
	.D(n_404),
	.Q(DPATH_RF_MEMORY_7__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_7__31_ (.CK(CTS_32),
	.D(n_403),
	.Q(DPATH_RF_MEMORY_7__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__0_ (.CK(CTS_19),
	.D(n_1037),
	.Q(DPATH_RF_MEMORY_8__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__1_ (.CK(CTS_50),
	.D(n_1040),
	.Q(DPATH_RF_MEMORY_8__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__2_ (.CK(CTS_11),
	.D(n_181),
	.Q(DPATH_RF_MEMORY_8__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__3_ (.CK(CTS_22),
	.D(n_1032),
	.Q(DPATH_RF_MEMORY_8__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__4_ (.CK(CTS_32),
	.D(n_1030),
	.Q(DPATH_RF_MEMORY_8__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__5_ (.CK(CTS_11),
	.D(n_1028),
	.Q(DPATH_RF_MEMORY_8__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__6_ (.CK(CTS_19),
	.D(n_1024),
	.Q(DPATH_RF_MEMORY_8__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__7_ (.CK(CTS_19),
	.D(n_1021),
	.Q(DPATH_RF_MEMORY_8__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__8_ (.CK(CTS_19),
	.D(n_1019),
	.Q(DPATH_RF_MEMORY_8__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__9_ (.CK(CTS_19),
	.D(n_1016),
	.Q(DPATH_RF_MEMORY_8__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__10_ (.CK(CTS_40),
	.D(n_1012),
	.Q(DPATH_RF_MEMORY_8__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__11_ (.CK(CTS_55),
	.D(n_1011),
	.Q(DPATH_RF_MEMORY_8__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__12_ (.CK(CTS_30),
	.D(n_1010),
	.Q(DPATH_RF_MEMORY_8__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__13_ (.CK(CTS_11),
	.D(n_1009),
	.Q(DPATH_RF_MEMORY_8__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__14_ (.CK(CTS_45),
	.D(n_1008),
	.Q(DPATH_RF_MEMORY_8__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__15_ (.CK(CTS_38),
	.D(n_1006),
	.Q(DPATH_RF_MEMORY_8__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__16_ (.CK(CTS_45),
	.D(n_1005),
	.Q(DPATH_RF_MEMORY_8__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__17_ (.CK(CTS_57),
	.D(n_1007),
	.Q(DPATH_RF_MEMORY_8__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__18_ (.CK(CTS_38),
	.D(n_1004),
	.Q(DPATH_RF_MEMORY_8__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__19_ (.CK(CTS_38),
	.D(n_1003),
	.Q(DPATH_RF_MEMORY_8__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__20_ (.CK(CTS_30),
	.D(n_1002),
	.Q(DPATH_RF_MEMORY_8__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__21_ (.CK(CTS_52),
	.D(n_1001),
	.Q(DPATH_RF_MEMORY_8__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__22_ (.CK(CTS_53),
	.D(n_1000),
	.Q(DPATH_RF_MEMORY_8__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__23_ (.CK(CTS_32),
	.D(n_999),
	.Q(DPATH_RF_MEMORY_8__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__24_ (.CK(CTS_55),
	.D(n_998),
	.Q(DPATH_RF_MEMORY_8__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__25_ (.CK(CTS_57),
	.D(n_997),
	.Q(DPATH_RF_MEMORY_8__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__26_ (.CK(CTS_43),
	.D(n_995),
	.Q(DPATH_RF_MEMORY_8__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__27_ (.CK(CTS_8),
	.D(n_992),
	.Q(DPATH_RF_MEMORY_8__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__28_ (.CK(CTS_4),
	.D(n_990),
	.Q(DPATH_RF_MEMORY_8__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__29_ (.CK(CTS_52),
	.D(n_989),
	.Q(DPATH_RF_MEMORY_8__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__30_ (.CK(CTS_56),
	.D(n_985),
	.Q(DPATH_RF_MEMORY_8__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_8__31_ (.CK(CTS_32),
	.D(n_979),
	.Q(DPATH_RF_MEMORY_8__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__0_ (.CK(CTS_18),
	.D(n_400),
	.Q(DPATH_RF_MEMORY_9__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__1_ (.CK(CTS_27),
	.D(n_401),
	.Q(DPATH_RF_MEMORY_9__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__2_ (.CK(CTS_27),
	.D(n_156),
	.Q(DPATH_RF_MEMORY_9__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__3_ (.CK(CTS_23),
	.D(n_399),
	.Q(DPATH_RF_MEMORY_9__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__4_ (.CK(CTS_32),
	.D(n_246),
	.Q(DPATH_RF_MEMORY_9__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__5_ (.CK(CTS_50),
	.D(n_398),
	.Q(DPATH_RF_MEMORY_9__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__6_ (.CK(CTS_60),
	.D(n_258),
	.Q(DPATH_RF_MEMORY_9__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__7_ (.CK(CTS_23),
	.D(n_397),
	.Q(DPATH_RF_MEMORY_9__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__8_ (.CK(CTS_18),
	.D(n_396),
	.Q(DPATH_RF_MEMORY_9__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__9_ (.CK(CTS_23),
	.D(n_395),
	.Q(DPATH_RF_MEMORY_9__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__10_ (.CK(CTS_40),
	.D(n_283),
	.Q(DPATH_RF_MEMORY_9__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__11_ (.CK(CTS_55),
	.D(n_394),
	.Q(DPATH_RF_MEMORY_9__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__12_ (.CK(CTS_4),
	.D(n_393),
	.Q(DPATH_RF_MEMORY_9__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__13_ (.CK(CTS_40),
	.D(n_392),
	.Q(DPATH_RF_MEMORY_9__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__14_ (.CK(CTS_46),
	.D(n_391),
	.Q(DPATH_RF_MEMORY_9__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__15_ (.CK(CTS_38),
	.D(n_387),
	.Q(DPATH_RF_MEMORY_9__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__16_ (.CK(CTS_46),
	.D(n_390),
	.Q(DPATH_RF_MEMORY_9__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__17_ (.CK(CTS_54),
	.D(n_388),
	.Q(DPATH_RF_MEMORY_9__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__18_ (.CK(CTS_54),
	.D(n_386),
	.Q(DPATH_RF_MEMORY_9__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__19_ (.CK(CTS_38),
	.D(n_385),
	.Q(DPATH_RF_MEMORY_9__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__20_ (.CK(CTS_21),
	.D(n_384),
	.Q(DPATH_RF_MEMORY_9__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__21_ (.CK(CTS_42),
	.D(n_383),
	.Q(DPATH_RF_MEMORY_9__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__22_ (.CK(CTS_42),
	.D(n_382),
	.Q(DPATH_RF_MEMORY_9__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__23_ (.CK(CTS_32),
	.D(n_381),
	.Q(DPATH_RF_MEMORY_9__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__24_ (.CK(CTS_47),
	.D(n_380),
	.Q(DPATH_RF_MEMORY_9__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__25_ (.CK(CTS_57),
	.D(n_379),
	.Q(DPATH_RF_MEMORY_9__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__26_ (.CK(CTS_3),
	.D(n_378),
	.Q(DPATH_RF_MEMORY_9__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__27_ (.CK(CTS_8),
	.D(n_377),
	.Q(DPATH_RF_MEMORY_9__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__28_ (.CK(CTS_17),
	.D(n_376),
	.Q(DPATH_RF_MEMORY_9__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__29_ (.CK(CTS_48),
	.D(n_375),
	.Q(DPATH_RF_MEMORY_9__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__30_ (.CK(CTS_47),
	.D(n_370),
	.Q(DPATH_RF_MEMORY_9__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_9__31_ (.CK(CTS_32),
	.D(n_373),
	.Q(DPATH_RF_MEMORY_9__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__0_ (.CK(CTS_18),
	.D(n_914),
	.Q(DPATH_RF_MEMORY_10__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__1_ (.CK(CTS_27),
	.D(n_917),
	.Q(DPATH_RF_MEMORY_10__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__2_ (.CK(CTS_27),
	.D(n_177),
	.Q(DPATH_RF_MEMORY_10__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__3_ (.CK(CTS_23),
	.D(n_909),
	.Q(DPATH_RF_MEMORY_10__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__4_ (.CK(CTS_32),
	.D(n_907),
	.Q(DPATH_RF_MEMORY_10__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__5_ (.CK(CTS_50),
	.D(n_906),
	.Q(DPATH_RF_MEMORY_10__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__6_ (.CK(CTS_60),
	.D(n_902),
	.Q(DPATH_RF_MEMORY_10__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__7_ (.CK(CTS_23),
	.D(n_900),
	.Q(DPATH_RF_MEMORY_10__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__8_ (.CK(CTS_18),
	.D(n_898),
	.Q(DPATH_RF_MEMORY_10__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__9_ (.CK(CTS_23),
	.D(n_895),
	.Q(DPATH_RF_MEMORY_10__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__10_ (.CK(CTS_40),
	.D(n_891),
	.Q(DPATH_RF_MEMORY_10__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__11_ (.CK(CTS_55),
	.D(n_890),
	.Q(DPATH_RF_MEMORY_10__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__12_ (.CK(CTS_4),
	.D(n_889),
	.Q(DPATH_RF_MEMORY_10__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__13_ (.CK(CTS_40),
	.D(n_888),
	.Q(DPATH_RF_MEMORY_10__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__14_ (.CK(CTS_46),
	.D(n_887),
	.Q(DPATH_RF_MEMORY_10__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__15_ (.CK(CTS_38),
	.D(n_886),
	.Q(DPATH_RF_MEMORY_10__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__16_ (.CK(CTS_46),
	.D(n_885),
	.Q(DPATH_RF_MEMORY_10__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__17_ (.CK(CTS_28),
	.D(n_884),
	.Q(DPATH_RF_MEMORY_10__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__18_ (.CK(CTS_54),
	.D(n_883),
	.Q(DPATH_RF_MEMORY_10__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__19_ (.CK(CTS_38),
	.D(n_882),
	.Q(DPATH_RF_MEMORY_10__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__20_ (.CK(CTS_29),
	.D(n_881),
	.Q(DPATH_RF_MEMORY_10__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__21_ (.CK(CTS_42),
	.D(n_880),
	.Q(DPATH_RF_MEMORY_10__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__22_ (.CK(CTS_42),
	.D(n_879),
	.Q(DPATH_RF_MEMORY_10__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__23_ (.CK(CTS_32),
	.D(n_878),
	.Q(DPATH_RF_MEMORY_10__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__24_ (.CK(CTS_53),
	.D(n_877),
	.Q(DPATH_RF_MEMORY_10__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__25_ (.CK(CTS_57),
	.D(n_876),
	.Q(DPATH_RF_MEMORY_10__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__26_ (.CK(CTS_3),
	.D(n_875),
	.Q(DPATH_RF_MEMORY_10__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__27_ (.CK(CTS_8),
	.D(n_874),
	.Q(DPATH_RF_MEMORY_10__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__28_ (.CK(CTS_17),
	.D(n_873),
	.Q(DPATH_RF_MEMORY_10__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__29_ (.CK(CTS_48),
	.D(n_872),
	.Q(DPATH_RF_MEMORY_10__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__30_ (.CK(CTS_45),
	.D(n_871),
	.Q(DPATH_RF_MEMORY_10__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_10__31_ (.CK(CTS_32),
	.D(n_870),
	.Q(DPATH_RF_MEMORY_10__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__0_ (.CK(CTS_22),
	.D(n_366),
	.Q(DPATH_RF_MEMORY_11__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__1_ (.CK(CTS_27),
	.D(n_365),
	.Q(DPATH_RF_MEMORY_11__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__2_ (.CK(CTS_27),
	.D(n_160),
	.Q(DPATH_RF_MEMORY_11__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__3_ (.CK(CTS_23),
	.D(n_363),
	.Q(DPATH_RF_MEMORY_11__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__4_ (.CK(CTS_32),
	.D(n_362),
	.Q(DPATH_RF_MEMORY_11__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__5_ (.CK(CTS_27),
	.D(n_361),
	.Q(DPATH_RF_MEMORY_11__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__6_ (.CK(CTS_60),
	.D(n_360),
	.Q(DPATH_RF_MEMORY_11__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__7_ (.CK(CTS_23),
	.D(n_359),
	.Q(DPATH_RF_MEMORY_11__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__8_ (.CK(CTS_23),
	.D(n_358),
	.Q(DPATH_RF_MEMORY_11__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__9_ (.CK(CTS_23),
	.D(n_357),
	.Q(DPATH_RF_MEMORY_11__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__10_ (.CK(CTS_40),
	.D(n_355),
	.Q(DPATH_RF_MEMORY_11__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__11_ (.CK(CTS_55),
	.D(n_353),
	.Q(DPATH_RF_MEMORY_11__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__12_ (.CK(CTS_59),
	.D(n_352),
	.Q(DPATH_RF_MEMORY_11__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__13_ (.CK(CTS_27),
	.D(n_351),
	.Q(DPATH_RF_MEMORY_11__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__14_ (.CK(CTS_48),
	.D(n_349),
	.Q(DPATH_RF_MEMORY_11__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__15_ (.CK(CTS_57),
	.D(n_348),
	.Q(DPATH_RF_MEMORY_11__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__16_ (.CK(CTS_47),
	.D(n_347),
	.Q(DPATH_RF_MEMORY_11__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__17_ (.CK(CTS_55),
	.D(n_346),
	.Q(DPATH_RF_MEMORY_11__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__18_ (.CK(CTS_54),
	.D(n_345),
	.Q(DPATH_RF_MEMORY_11__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__19_ (.CK(CTS_38),
	.D(n_344),
	.Q(DPATH_RF_MEMORY_11__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__20_ (.CK(CTS_21),
	.D(n_343),
	.Q(DPATH_RF_MEMORY_11__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__21_ (.CK(CTS_42),
	.D(n_342),
	.Q(DPATH_RF_MEMORY_11__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__22_ (.CK(CTS_48),
	.D(n_341),
	.Q(DPATH_RF_MEMORY_11__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__23_ (.CK(CTS_8),
	.D(n_339),
	.Q(DPATH_RF_MEMORY_11__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__24_ (.CK(CTS_47),
	.D(n_338),
	.Q(DPATH_RF_MEMORY_11__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__25_ (.CK(CTS_57),
	.D(n_337),
	.Q(DPATH_RF_MEMORY_11__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__26_ (.CK(CTS_3),
	.D(n_336),
	.Q(DPATH_RF_MEMORY_11__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__27_ (.CK(CTS_26),
	.D(n_334),
	.Q(DPATH_RF_MEMORY_11__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__28_ (.CK(CTS_17),
	.D(n_332),
	.Q(DPATH_RF_MEMORY_11__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__29_ (.CK(CTS_48),
	.D(n_331),
	.Q(DPATH_RF_MEMORY_11__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__30_ (.CK(CTS_47),
	.D(n_330),
	.Q(DPATH_RF_MEMORY_11__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_11__31_ (.CK(CTS_32),
	.D(n_329),
	.Q(DPATH_RF_MEMORY_11__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__0_ (.CK(CTS_18),
	.D(n_869),
	.Q(DPATH_RF_MEMORY_12__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__1_ (.CK(CTS_27),
	.D(n_868),
	.Q(DPATH_RF_MEMORY_12__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__2_ (.CK(CTS_50),
	.D(n_176),
	.Q(DPATH_RF_MEMORY_12__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__3_ (.CK(CTS_22),
	.D(n_867),
	.Q(DPATH_RF_MEMORY_12__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__4_ (.CK(CTS_32),
	.D(n_866),
	.Q(DPATH_RF_MEMORY_12__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__5_ (.CK(CTS_27),
	.D(n_865),
	.Q(DPATH_RF_MEMORY_12__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__6_ (.CK(CTS_60),
	.D(n_864),
	.Q(DPATH_RF_MEMORY_12__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__7_ (.CK(CTS_22),
	.D(n_863),
	.Q(DPATH_RF_MEMORY_12__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__8_ (.CK(CTS_22),
	.D(n_862),
	.Q(DPATH_RF_MEMORY_12__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__9_ (.CK(CTS_23),
	.D(n_861),
	.Q(DPATH_RF_MEMORY_12__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__10_ (.CK(CTS_40),
	.D(n_860),
	.Q(DPATH_RF_MEMORY_12__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__11_ (.CK(CTS_55),
	.D(n_859),
	.Q(DPATH_RF_MEMORY_12__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__12_ (.CK(CTS_59),
	.D(n_858),
	.Q(DPATH_RF_MEMORY_12__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__13_ (.CK(CTS_40),
	.D(n_857),
	.Q(DPATH_RF_MEMORY_12__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__14_ (.CK(CTS_48),
	.D(n_856),
	.Q(DPATH_RF_MEMORY_12__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__15_ (.CK(CTS_57),
	.D(n_855),
	.Q(DPATH_RF_MEMORY_12__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__16_ (.CK(CTS_46),
	.D(n_854),
	.Q(DPATH_RF_MEMORY_12__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__17_ (.CK(CTS_28),
	.D(n_853),
	.Q(DPATH_RF_MEMORY_12__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__18_ (.CK(CTS_54),
	.D(n_852),
	.Q(DPATH_RF_MEMORY_12__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__19_ (.CK(CTS_38),
	.D(n_851),
	.Q(DPATH_RF_MEMORY_12__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__20_ (.CK(CTS_21),
	.D(n_850),
	.Q(DPATH_RF_MEMORY_12__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__21_ (.CK(CTS_42),
	.D(n_849),
	.Q(DPATH_RF_MEMORY_12__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__22_ (.CK(CTS_48),
	.D(n_848),
	.Q(DPATH_RF_MEMORY_12__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__23_ (.CK(CTS_8),
	.D(n_847),
	.Q(DPATH_RF_MEMORY_12__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__24_ (.CK(CTS_53),
	.D(n_846),
	.Q(DPATH_RF_MEMORY_12__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__25_ (.CK(CTS_57),
	.D(n_845),
	.Q(DPATH_RF_MEMORY_12__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__26_ (.CK(CTS_3),
	.D(n_844),
	.Q(DPATH_RF_MEMORY_12__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__27_ (.CK(CTS_8),
	.D(n_843),
	.Q(DPATH_RF_MEMORY_12__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__28_ (.CK(CTS_17),
	.D(n_842),
	.Q(DPATH_RF_MEMORY_12__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__29_ (.CK(CTS_48),
	.D(n_841),
	.Q(DPATH_RF_MEMORY_12__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__30_ (.CK(CTS_45),
	.D(n_840),
	.Q(DPATH_RF_MEMORY_12__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_12__31_ (.CK(CTS_32),
	.D(n_839),
	.Q(DPATH_RF_MEMORY_12__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__0_ (.CK(CTS_18),
	.D(n_521),
	.Q(DPATH_RF_MEMORY_13__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__1_ (.CK(CTS_27),
	.D(n_520),
	.Q(DPATH_RF_MEMORY_13__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__2_ (.CK(CTS_27),
	.D(n_166),
	.Q(DPATH_RF_MEMORY_13__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__3_ (.CK(CTS_23),
	.D(n_519),
	.Q(DPATH_RF_MEMORY_13__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__4_ (.CK(CTS_17),
	.D(n_518),
	.Q(DPATH_RF_MEMORY_13__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__5_ (.CK(CTS_50),
	.D(n_517),
	.Q(DPATH_RF_MEMORY_13__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__6_ (.CK(CTS_60),
	.D(n_516),
	.Q(DPATH_RF_MEMORY_13__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__7_ (.CK(CTS_23),
	.D(n_515),
	.Q(DPATH_RF_MEMORY_13__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__8_ (.CK(CTS_18),
	.D(n_514),
	.Q(DPATH_RF_MEMORY_13__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__9_ (.CK(CTS_23),
	.D(n_513),
	.Q(DPATH_RF_MEMORY_13__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__10_ (.CK(CTS_27),
	.D(n_512),
	.Q(DPATH_RF_MEMORY_13__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__11_ (.CK(CTS_54),
	.D(n_511),
	.Q(DPATH_RF_MEMORY_13__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__12_ (.CK(CTS_3),
	.D(n_510),
	.Q(DPATH_RF_MEMORY_13__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__13_ (.CK(CTS_40),
	.D(n_509),
	.Q(DPATH_RF_MEMORY_13__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__14_ (.CK(CTS_48),
	.D(n_506),
	.Q(DPATH_RF_MEMORY_13__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__15_ (.CK(CTS_54),
	.D(n_508),
	.Q(DPATH_RF_MEMORY_13__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__16_ (.CK(CTS_46),
	.D(n_507),
	.Q(DPATH_RF_MEMORY_13__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__17_ (.CK(CTS_54),
	.D(n_505),
	.Q(DPATH_RF_MEMORY_13__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__18_ (.CK(CTS_54),
	.D(n_504),
	.Q(DPATH_RF_MEMORY_13__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__19_ (.CK(CTS_26),
	.D(n_503),
	.Q(DPATH_RF_MEMORY_13__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__20_ (.CK(CTS_13),
	.D(n_502),
	.Q(DPATH_RF_MEMORY_13__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__21_ (.CK(CTS_48),
	.D(n_501),
	.Q(DPATH_RF_MEMORY_13__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__22_ (.CK(CTS_48),
	.D(n_500),
	.Q(DPATH_RF_MEMORY_13__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__23_ (.CK(CTS_8),
	.D(n_499),
	.Q(DPATH_RF_MEMORY_13__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__24_ (.CK(CTS_47),
	.D(n_498),
	.Q(DPATH_RF_MEMORY_13__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__25_ (.CK(CTS_57),
	.D(n_497),
	.Q(DPATH_RF_MEMORY_13__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__26_ (.CK(CTS_3),
	.D(n_496),
	.Q(DPATH_RF_MEMORY_13__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__27_ (.CK(CTS_26),
	.D(n_495),
	.Q(DPATH_RF_MEMORY_13__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__28_ (.CK(CTS_29),
	.D(n_494),
	.Q(DPATH_RF_MEMORY_13__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__29_ (.CK(CTS_48),
	.D(n_493),
	.Q(DPATH_RF_MEMORY_13__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__30_ (.CK(CTS_47),
	.D(n_492),
	.Q(DPATH_RF_MEMORY_13__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_13__31_ (.CK(CTS_17),
	.D(n_491),
	.Q(DPATH_RF_MEMORY_13__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__0_ (.CK(CTS_18),
	.D(n_838),
	.Q(DPATH_RF_MEMORY_14__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__1_ (.CK(CTS_60),
	.D(n_837),
	.Q(DPATH_RF_MEMORY_14__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__2_ (.CK(CTS_27),
	.D(n_175),
	.Q(DPATH_RF_MEMORY_14__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__3_ (.CK(CTS_23),
	.D(n_836),
	.Q(DPATH_RF_MEMORY_14__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__4_ (.CK(CTS_17),
	.D(n_835),
	.Q(DPATH_RF_MEMORY_14__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__5_ (.CK(CTS_41),
	.D(n_834),
	.Q(DPATH_RF_MEMORY_14__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__6_ (.CK(CTS_60),
	.D(n_833),
	.Q(DPATH_RF_MEMORY_14__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__7_ (.CK(CTS_23),
	.D(n_832),
	.Q(DPATH_RF_MEMORY_14__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__8_ (.CK(CTS_18),
	.D(n_831),
	.Q(DPATH_RF_MEMORY_14__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__9_ (.CK(CTS_23),
	.D(n_830),
	.Q(DPATH_RF_MEMORY_14__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__10_ (.CK(CTS_27),
	.D(n_829),
	.Q(DPATH_RF_MEMORY_14__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__11_ (.CK(CTS_55),
	.D(n_828),
	.Q(DPATH_RF_MEMORY_14__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__12_ (.CK(CTS_3),
	.D(n_827),
	.Q(DPATH_RF_MEMORY_14__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__13_ (.CK(CTS_40),
	.D(n_826),
	.Q(DPATH_RF_MEMORY_14__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__14_ (.CK(CTS_48),
	.D(n_825),
	.Q(DPATH_RF_MEMORY_14__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__15_ (.CK(CTS_28),
	.D(n_824),
	.Q(DPATH_RF_MEMORY_14__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__16_ (.CK(CTS_46),
	.D(n_823),
	.Q(DPATH_RF_MEMORY_14__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__17_ (.CK(CTS_55),
	.D(n_822),
	.Q(DPATH_RF_MEMORY_14__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__18_ (.CK(CTS_54),
	.D(n_821),
	.Q(DPATH_RF_MEMORY_14__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__19_ (.CK(CTS_28),
	.D(n_820),
	.Q(DPATH_RF_MEMORY_14__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__20_ (.CK(CTS_21),
	.D(n_819),
	.Q(DPATH_RF_MEMORY_14__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__21_ (.CK(CTS_42),
	.D(n_818),
	.Q(DPATH_RF_MEMORY_14__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__22_ (.CK(CTS_48),
	.D(n_817),
	.Q(DPATH_RF_MEMORY_14__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__23_ (.CK(CTS_21),
	.D(n_816),
	.Q(DPATH_RF_MEMORY_14__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__24_ (.CK(CTS_56),
	.D(n_815),
	.Q(DPATH_RF_MEMORY_14__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__25_ (.CK(CTS_54),
	.D(n_814),
	.Q(DPATH_RF_MEMORY_14__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__26_ (.CK(CTS_9),
	.D(n_813),
	.Q(DPATH_RF_MEMORY_14__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__27_ (.CK(CTS_26),
	.D(n_812),
	.Q(DPATH_RF_MEMORY_14__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__28_ (.CK(CTS_29),
	.D(n_811),
	.Q(DPATH_RF_MEMORY_14__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__29_ (.CK(CTS_48),
	.D(n_810),
	.Q(DPATH_RF_MEMORY_14__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__30_ (.CK(CTS_47),
	.D(n_809),
	.Q(DPATH_RF_MEMORY_14__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_14__31_ (.CK(CTS_17),
	.D(n_808),
	.Q(DPATH_RF_MEMORY_14__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__0_ (.CK(CTS_18),
	.D(n_312),
	.Q(DPATH_RF_MEMORY_15__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__1_ (.CK(CTS_27),
	.D(n_311),
	.Q(DPATH_RF_MEMORY_15__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__2_ (.CK(CTS_27),
	.D(n_159),
	.Q(DPATH_RF_MEMORY_15__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__3_ (.CK(CTS_22),
	.D(n_310),
	.Q(DPATH_RF_MEMORY_15__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__4_ (.CK(CTS_17),
	.D(n_309),
	.Q(DPATH_RF_MEMORY_15__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__5_ (.CK(CTS_50),
	.D(n_308),
	.Q(DPATH_RF_MEMORY_15__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__6_ (.CK(CTS_60),
	.D(n_307),
	.Q(DPATH_RF_MEMORY_15__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__7_ (.CK(CTS_23),
	.D(n_306),
	.Q(DPATH_RF_MEMORY_15__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__8_ (.CK(CTS_22),
	.D(n_305),
	.Q(DPATH_RF_MEMORY_15__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__9_ (.CK(CTS_23),
	.D(n_304),
	.Q(DPATH_RF_MEMORY_15__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__10_ (.CK(CTS_27),
	.D(n_303),
	.Q(DPATH_RF_MEMORY_15__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__11_ (.CK(CTS_56),
	.D(n_302),
	.Q(DPATH_RF_MEMORY_15__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__12_ (.CK(CTS_4),
	.D(n_301),
	.Q(DPATH_RF_MEMORY_15__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__13_ (.CK(CTS_50),
	.D(n_300),
	.Q(DPATH_RF_MEMORY_15__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__14_ (.CK(CTS_48),
	.D(n_299),
	.Q(DPATH_RF_MEMORY_15__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__15_ (.CK(CTS_54),
	.D(n_298),
	.Q(DPATH_RF_MEMORY_15__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__16_ (.CK(CTS_48),
	.D(n_297),
	.Q(DPATH_RF_MEMORY_15__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__17_ (.CK(CTS_54),
	.D(n_296),
	.Q(DPATH_RF_MEMORY_15__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__18_ (.CK(CTS_54),
	.D(n_295),
	.Q(DPATH_RF_MEMORY_15__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__19_ (.CK(CTS_28),
	.D(n_294),
	.Q(DPATH_RF_MEMORY_15__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__20_ (.CK(CTS_29),
	.D(n_293),
	.Q(DPATH_RF_MEMORY_15__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__21_ (.CK(CTS_48),
	.D(n_292),
	.Q(DPATH_RF_MEMORY_15__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__22_ (.CK(CTS_48),
	.D(n_291),
	.Q(DPATH_RF_MEMORY_15__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__23_ (.CK(CTS_21),
	.D(n_290),
	.Q(DPATH_RF_MEMORY_15__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__24_ (.CK(CTS_47),
	.D(n_289),
	.Q(DPATH_RF_MEMORY_15__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__25_ (.CK(CTS_54),
	.D(n_288),
	.Q(DPATH_RF_MEMORY_15__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__26_ (.CK(CTS_3),
	.D(n_287),
	.Q(DPATH_RF_MEMORY_15__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__27_ (.CK(CTS_8),
	.D(n_286),
	.Q(DPATH_RF_MEMORY_15__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__28_ (.CK(CTS_17),
	.D(n_285),
	.Q(DPATH_RF_MEMORY_15__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__29_ (.CK(CTS_48),
	.D(n_284),
	.Q(DPATH_RF_MEMORY_15__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__30_ (.CK(CTS_47),
	.D(n_282),
	.Q(DPATH_RF_MEMORY_15__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_15__31_ (.CK(CTS_21),
	.D(n_281),
	.Q(DPATH_RF_MEMORY_15__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__0_ (.CK(CTS_18),
	.D(n_807),
	.Q(DPATH_RF_MEMORY_16__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__1_ (.CK(CTS_27),
	.D(n_806),
	.Q(DPATH_RF_MEMORY_16__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__2_ (.CK(CTS_27),
	.D(n_174),
	.Q(DPATH_RF_MEMORY_16__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__3_ (.CK(CTS_22),
	.D(n_805),
	.Q(DPATH_RF_MEMORY_16__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__4_ (.CK(CTS_17),
	.D(n_804),
	.Q(DPATH_RF_MEMORY_16__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__5_ (.CK(CTS_50),
	.D(n_803),
	.Q(DPATH_RF_MEMORY_16__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__6_ (.CK(CTS_60),
	.D(n_802),
	.Q(DPATH_RF_MEMORY_16__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__7_ (.CK(CTS_23),
	.D(n_801),
	.Q(DPATH_RF_MEMORY_16__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__8_ (.CK(CTS_18),
	.D(n_800),
	.Q(DPATH_RF_MEMORY_16__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__9_ (.CK(CTS_23),
	.D(n_799),
	.Q(DPATH_RF_MEMORY_16__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__10_ (.CK(CTS_27),
	.D(n_798),
	.Q(DPATH_RF_MEMORY_16__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__11_ (.CK(CTS_55),
	.D(n_797),
	.Q(DPATH_RF_MEMORY_16__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__12_ (.CK(CTS_4),
	.D(n_796),
	.Q(DPATH_RF_MEMORY_16__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__13_ (.CK(CTS_50),
	.D(n_795),
	.Q(DPATH_RF_MEMORY_16__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__14_ (.CK(CTS_46),
	.D(n_794),
	.Q(DPATH_RF_MEMORY_16__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__15_ (.CK(CTS_28),
	.D(n_793),
	.Q(DPATH_RF_MEMORY_16__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__16_ (.CK(CTS_46),
	.D(n_792),
	.Q(DPATH_RF_MEMORY_16__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__17_ (.CK(CTS_55),
	.D(n_791),
	.Q(DPATH_RF_MEMORY_16__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__18_ (.CK(CTS_54),
	.D(n_790),
	.Q(DPATH_RF_MEMORY_16__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__19_ (.CK(CTS_28),
	.D(n_789),
	.Q(DPATH_RF_MEMORY_16__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__20_ (.CK(CTS_29),
	.D(n_788),
	.Q(DPATH_RF_MEMORY_16__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__21_ (.CK(CTS_48),
	.D(n_787),
	.Q(DPATH_RF_MEMORY_16__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__22_ (.CK(CTS_48),
	.D(n_786),
	.Q(DPATH_RF_MEMORY_16__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__23_ (.CK(CTS_29),
	.D(n_785),
	.Q(DPATH_RF_MEMORY_16__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__24_ (.CK(CTS_47),
	.D(n_784),
	.Q(DPATH_RF_MEMORY_16__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__25_ (.CK(CTS_54),
	.D(n_783),
	.Q(DPATH_RF_MEMORY_16__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__26_ (.CK(CTS_3),
	.D(n_782),
	.Q(DPATH_RF_MEMORY_16__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__27_ (.CK(CTS_21),
	.D(n_781),
	.Q(DPATH_RF_MEMORY_16__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__28_ (.CK(CTS_17),
	.D(n_780),
	.Q(DPATH_RF_MEMORY_16__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__29_ (.CK(CTS_48),
	.D(n_779),
	.Q(DPATH_RF_MEMORY_16__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__30_ (.CK(CTS_47),
	.D(n_778),
	.Q(DPATH_RF_MEMORY_16__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_16__31_ (.CK(CTS_21),
	.D(n_777),
	.Q(DPATH_RF_MEMORY_16__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__0_ (.CK(CTS_15),
	.D(n_269),
	.Q(DPATH_RF_MEMORY_17__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__1_ (.CK(CTS_16),
	.D(n_267),
	.Q(DPATH_RF_MEMORY_17__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__2_ (.CK(CTS_41),
	.D(n_157),
	.Q(DPATH_RF_MEMORY_17__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__3_ (.CK(CTS_22),
	.D(n_265),
	.Q(DPATH_RF_MEMORY_17__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__4_ (.CK(CTS_29),
	.D(n_264),
	.Q(DPATH_RF_MEMORY_17__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__5_ (.CK(CTS_16),
	.D(n_263),
	.Q(DPATH_RF_MEMORY_17__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__6_ (.CK(CTS_15),
	.D(n_261),
	.Q(DPATH_RF_MEMORY_17__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__7_ (.CK(CTS_22),
	.D(n_259),
	.Q(DPATH_RF_MEMORY_17__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__8_ (.CK(CTS_22),
	.D(n_256),
	.Q(DPATH_RF_MEMORY_17__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__9_ (.CK(CTS_22),
	.D(n_255),
	.Q(DPATH_RF_MEMORY_17__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__10_ (.CK(CTS_41),
	.D(n_254),
	.Q(DPATH_RF_MEMORY_17__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__11_ (.CK(CTS_52),
	.D(n_252),
	.Q(DPATH_RF_MEMORY_17__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__12_ (.CK(CTS_59),
	.D(n_250),
	.Q(DPATH_RF_MEMORY_17__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__13_ (.CK(CTS_41),
	.D(n_249),
	.Q(DPATH_RF_MEMORY_17__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__14_ (.CK(CTS_42),
	.D(n_248),
	.Q(DPATH_RF_MEMORY_17__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__15_ (.CK(CTS_26),
	.D(n_247),
	.Q(DPATH_RF_MEMORY_17__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__16_ (.CK(CTS_45),
	.D(n_245),
	.Q(DPATH_RF_MEMORY_17__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__17_ (.CK(CTS_28),
	.D(n_243),
	.Q(DPATH_RF_MEMORY_17__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__18_ (.CK(CTS_28),
	.D(n_241),
	.Q(DPATH_RF_MEMORY_17__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__19_ (.CK(CTS_26),
	.D(n_239),
	.Q(DPATH_RF_MEMORY_17__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__20_ (.CK(CTS_21),
	.D(n_238),
	.Q(DPATH_RF_MEMORY_17__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__21_ (.CK(CTS_42),
	.D(n_237),
	.Q(DPATH_RF_MEMORY_17__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__22_ (.CK(CTS_42),
	.D(n_235),
	.Q(DPATH_RF_MEMORY_17__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__23_ (.CK(CTS_8),
	.D(n_233),
	.Q(DPATH_RF_MEMORY_17__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__24_ (.CK(CTS_51),
	.D(n_231),
	.Q(DPATH_RF_MEMORY_17__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__25_ (.CK(CTS_28),
	.D(n_230),
	.Q(DPATH_RF_MEMORY_17__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__26_ (.CK(CTS_3),
	.D(n_229),
	.Q(DPATH_RF_MEMORY_17__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__27_ (.CK(CTS_8),
	.D(n_227),
	.Q(DPATH_RF_MEMORY_17__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__28_ (.CK(CTS_59),
	.D(n_226),
	.Q(DPATH_RF_MEMORY_17__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__29_ (.CK(CTS_45),
	.D(n_224),
	.Q(DPATH_RF_MEMORY_17__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__30_ (.CK(CTS_51),
	.D(n_222),
	.Q(DPATH_RF_MEMORY_17__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_17__31_ (.CK(CTS_32),
	.D(n_221),
	.Q(DPATH_RF_MEMORY_17__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__0_ (.CK(CTS_19),
	.D(n_776),
	.Q(DPATH_RF_MEMORY_18__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__1_ (.CK(CTS_16),
	.D(n_775),
	.Q(DPATH_RF_MEMORY_18__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__2_ (.CK(CTS_40),
	.D(n_173),
	.Q(DPATH_RF_MEMORY_18__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__3_ (.CK(CTS_22),
	.D(n_774),
	.Q(DPATH_RF_MEMORY_18__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__4_ (.CK(CTS_32),
	.D(n_773),
	.Q(DPATH_RF_MEMORY_18__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__5_ (.CK(CTS_50),
	.D(n_772),
	.Q(DPATH_RF_MEMORY_18__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__6_ (.CK(CTS_15),
	.D(n_771),
	.Q(DPATH_RF_MEMORY_18__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__7_ (.CK(CTS_22),
	.D(n_770),
	.Q(DPATH_RF_MEMORY_18__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__8_ (.CK(CTS_22),
	.D(n_768),
	.Q(DPATH_RF_MEMORY_18__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__9_ (.CK(CTS_19),
	.D(n_767),
	.Q(DPATH_RF_MEMORY_18__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__10_ (.CK(CTS_41),
	.D(n_766),
	.Q(DPATH_RF_MEMORY_18__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__11_ (.CK(CTS_52),
	.D(n_765),
	.Q(DPATH_RF_MEMORY_18__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__12_ (.CK(CTS_59),
	.D(n_764),
	.Q(DPATH_RF_MEMORY_18__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__13_ (.CK(CTS_40),
	.D(n_763),
	.Q(DPATH_RF_MEMORY_18__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__14_ (.CK(CTS_45),
	.D(n_762),
	.Q(DPATH_RF_MEMORY_18__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__15_ (.CK(CTS_38),
	.D(n_761),
	.Q(DPATH_RF_MEMORY_18__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__16_ (.CK(CTS_45),
	.D(n_759),
	.Q(DPATH_RF_MEMORY_18__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__17_ (.CK(CTS_28),
	.D(n_758),
	.Q(DPATH_RF_MEMORY_18__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__18_ (.CK(CTS_28),
	.D(n_755),
	.Q(DPATH_RF_MEMORY_18__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__19_ (.CK(CTS_8),
	.D(n_754),
	.Q(DPATH_RF_MEMORY_18__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__20_ (.CK(CTS_21),
	.D(n_753),
	.Q(DPATH_RF_MEMORY_18__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__21_ (.CK(CTS_52),
	.D(n_752),
	.Q(DPATH_RF_MEMORY_18__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__22_ (.CK(CTS_46),
	.D(n_749),
	.Q(DPATH_RF_MEMORY_18__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__23_ (.CK(CTS_32),
	.D(n_748),
	.Q(DPATH_RF_MEMORY_18__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__24_ (.CK(CTS_45),
	.D(n_746),
	.Q(DPATH_RF_MEMORY_18__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__25_ (.CK(CTS_8),
	.D(n_745),
	.Q(DPATH_RF_MEMORY_18__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__26_ (.CK(CTS_9),
	.D(n_743),
	.Q(DPATH_RF_MEMORY_18__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__27_ (.CK(CTS_8),
	.D(n_742),
	.Q(DPATH_RF_MEMORY_18__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__28_ (.CK(CTS_59),
	.D(n_741),
	.Q(DPATH_RF_MEMORY_18__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__29_ (.CK(CTS_51),
	.D(n_739),
	.Q(DPATH_RF_MEMORY_18__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__30_ (.CK(CTS_53),
	.D(n_737),
	.Q(DPATH_RF_MEMORY_18__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_18__31_ (.CK(CTS_32),
	.D(n_736),
	.Q(DPATH_RF_MEMORY_18__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__0_ (.CK(CTS_18),
	.D(n_216),
	.Q(DPATH_RF_MEMORY_19__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__1_ (.CK(CTS_16),
	.D(n_215),
	.Q(DPATH_RF_MEMORY_19__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__2_ (.CK(CTS_41),
	.D(n_155),
	.Q(DPATH_RF_MEMORY_19__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__3_ (.CK(CTS_1),
	.D(n_214),
	.Q(DPATH_RF_MEMORY_19__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__4_ (.CK(CTS_29),
	.D(n_213),
	.Q(DPATH_RF_MEMORY_19__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__5_ (.CK(CTS_41),
	.D(n_212),
	.Q(DPATH_RF_MEMORY_19__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__6_ (.CK(CTS_15),
	.D(n_211),
	.Q(DPATH_RF_MEMORY_19__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__7_ (.CK(CTS_1),
	.D(n_210),
	.Q(DPATH_RF_MEMORY_19__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__8_ (.CK(CTS_1),
	.D(n_209),
	.Q(DPATH_RF_MEMORY_19__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__9_ (.CK(CTS_1),
	.D(n_208),
	.Q(DPATH_RF_MEMORY_19__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__10_ (.CK(CTS_41),
	.D(n_207),
	.Q(DPATH_RF_MEMORY_19__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__11_ (.CK(CTS_52),
	.D(n_206),
	.Q(DPATH_RF_MEMORY_19__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__12_ (.CK(CTS_3),
	.D(n_205),
	.Q(DPATH_RF_MEMORY_19__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__13_ (.CK(CTS_41),
	.D(n_204),
	.Q(DPATH_RF_MEMORY_19__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__14_ (.CK(CTS_46),
	.D(n_203),
	.Q(DPATH_RF_MEMORY_19__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__15_ (.CK(CTS_26),
	.D(n_202),
	.Q(DPATH_RF_MEMORY_19__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__16_ (.CK(CTS_45),
	.D(n_201),
	.Q(DPATH_RF_MEMORY_19__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__17_ (.CK(CTS_28),
	.D(n_200),
	.Q(DPATH_RF_MEMORY_19__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__18_ (.CK(CTS_28),
	.D(n_199),
	.Q(DPATH_RF_MEMORY_19__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__19_ (.CK(CTS_26),
	.D(n_198),
	.Q(DPATH_RF_MEMORY_19__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__20_ (.CK(CTS_13),
	.D(n_197),
	.Q(DPATH_RF_MEMORY_19__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__21_ (.CK(CTS_42),
	.D(n_196),
	.Q(DPATH_RF_MEMORY_19__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__22_ (.CK(CTS_45),
	.D(n_195),
	.Q(DPATH_RF_MEMORY_19__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__23_ (.CK(CTS_21),
	.D(n_194),
	.Q(DPATH_RF_MEMORY_19__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__24_ (.CK(CTS_45),
	.D(n_193),
	.Q(DPATH_RF_MEMORY_19__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__25_ (.CK(CTS_28),
	.D(n_192),
	.Q(DPATH_RF_MEMORY_19__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__26_ (.CK(CTS_9),
	.D(n_191),
	.Q(DPATH_RF_MEMORY_19__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__27_ (.CK(CTS_21),
	.D(n_190),
	.Q(DPATH_RF_MEMORY_19__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__28_ (.CK(CTS_29),
	.D(n_189),
	.Q(DPATH_RF_MEMORY_19__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__29_ (.CK(CTS_45),
	.D(n_188),
	.Q(DPATH_RF_MEMORY_19__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__30_ (.CK(CTS_53),
	.D(n_187),
	.Q(DPATH_RF_MEMORY_19__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_19__31_ (.CK(CTS_17),
	.D(n_186),
	.Q(DPATH_RF_MEMORY_19__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__0_ (.CK(CTS_1),
	.D(n_717),
	.Q(DPATH_RF_MEMORY_20__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__1_ (.CK(CTS_16),
	.D(n_716),
	.Q(DPATH_RF_MEMORY_20__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__2_ (.CK(CTS_41),
	.D(n_171),
	.Q(DPATH_RF_MEMORY_20__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__3_ (.CK(CTS_5),
	.D(n_714),
	.Q(DPATH_RF_MEMORY_20__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__4_ (.CK(CTS_17),
	.D(n_713),
	.Q(DPATH_RF_MEMORY_20__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__5_ (.CK(CTS_16),
	.D(n_711),
	.Q(DPATH_RF_MEMORY_20__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__6_ (.CK(CTS_16),
	.D(n_709),
	.Q(DPATH_RF_MEMORY_20__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__7_ (.CK(CTS_1),
	.D(n_707),
	.Q(DPATH_RF_MEMORY_20__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__8_ (.CK(CTS_1),
	.D(n_706),
	.Q(DPATH_RF_MEMORY_20__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__9_ (.CK(CTS_1),
	.D(n_705),
	.Q(DPATH_RF_MEMORY_20__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__10_ (.CK(CTS_41),
	.D(n_704),
	.Q(DPATH_RF_MEMORY_20__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__11_ (.CK(CTS_52),
	.D(n_702),
	.Q(DPATH_RF_MEMORY_20__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__12_ (.CK(CTS_59),
	.D(n_701),
	.Q(DPATH_RF_MEMORY_20__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__13_ (.CK(CTS_41),
	.D(n_700),
	.Q(DPATH_RF_MEMORY_20__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__14_ (.CK(CTS_45),
	.D(n_699),
	.Q(DPATH_RF_MEMORY_20__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__15_ (.CK(CTS_28),
	.D(n_698),
	.Q(DPATH_RF_MEMORY_20__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__16_ (.CK(CTS_45),
	.D(n_697),
	.Q(DPATH_RF_MEMORY_20__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__17_ (.CK(CTS_28),
	.D(n_696),
	.Q(DPATH_RF_MEMORY_20__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__18_ (.CK(CTS_13),
	.D(n_695),
	.Q(DPATH_RF_MEMORY_20__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__19_ (.CK(CTS_13),
	.D(n_694),
	.Q(DPATH_RF_MEMORY_20__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__20_ (.CK(CTS_13),
	.D(n_693),
	.Q(DPATH_RF_MEMORY_20__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__21_ (.CK(CTS_42),
	.D(n_692),
	.Q(DPATH_RF_MEMORY_20__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__22_ (.CK(CTS_42),
	.D(n_691),
	.Q(DPATH_RF_MEMORY_20__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__23_ (.CK(CTS_21),
	.D(n_690),
	.Q(DPATH_RF_MEMORY_20__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__24_ (.CK(CTS_45),
	.D(n_689),
	.Q(DPATH_RF_MEMORY_20__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__25_ (.CK(CTS_13),
	.D(n_688),
	.Q(DPATH_RF_MEMORY_20__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__26_ (.CK(CTS_3),
	.D(n_687),
	.Q(DPATH_RF_MEMORY_20__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__27_ (.CK(CTS_13),
	.D(n_686),
	.Q(DPATH_RF_MEMORY_20__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__28_ (.CK(CTS_29),
	.D(n_685),
	.Q(DPATH_RF_MEMORY_20__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__29_ (.CK(CTS_46),
	.D(n_684),
	.Q(DPATH_RF_MEMORY_20__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__30_ (.CK(CTS_53),
	.D(n_683),
	.Q(DPATH_RF_MEMORY_20__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_20__31_ (.CK(CTS_29),
	.D(n_682),
	.Q(DPATH_RF_MEMORY_20__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__0_ (.CK(CTS_18),
	.D(n_479),
	.Q(DPATH_RF_MEMORY_21__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__1_ (.CK(CTS_16),
	.D(n_478),
	.Q(DPATH_RF_MEMORY_21__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__2_ (.CK(CTS_41),
	.D(n_164),
	.Q(DPATH_RF_MEMORY_21__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__3_ (.CK(CTS_1),
	.D(n_476),
	.Q(DPATH_RF_MEMORY_21__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__4_ (.CK(CTS_29),
	.D(n_475),
	.Q(DPATH_RF_MEMORY_21__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__5_ (.CK(CTS_16),
	.D(n_473),
	.Q(DPATH_RF_MEMORY_21__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__6_ (.CK(CTS_15),
	.D(n_471),
	.Q(DPATH_RF_MEMORY_21__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__7_ (.CK(CTS_1),
	.D(n_469),
	.Q(DPATH_RF_MEMORY_21__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__8_ (.CK(CTS_18),
	.D(n_468),
	.Q(DPATH_RF_MEMORY_21__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__9_ (.CK(CTS_19),
	.D(n_467),
	.Q(DPATH_RF_MEMORY_21__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__10_ (.CK(CTS_40),
	.D(n_465),
	.Q(DPATH_RF_MEMORY_21__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__11_ (.CK(CTS_52),
	.D(n_556),
	.Q(DPATH_RF_MEMORY_21__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__12_ (.CK(CTS_9),
	.D(n_555),
	.Q(DPATH_RF_MEMORY_21__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__13_ (.CK(CTS_41),
	.D(n_554),
	.Q(DPATH_RF_MEMORY_21__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__14_ (.CK(CTS_45),
	.D(n_553),
	.Q(DPATH_RF_MEMORY_21__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__15_ (.CK(CTS_26),
	.D(n_552),
	.Q(DPATH_RF_MEMORY_21__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__16_ (.CK(CTS_51),
	.D(n_550),
	.Q(DPATH_RF_MEMORY_21__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__17_ (.CK(CTS_28),
	.D(n_548),
	.Q(DPATH_RF_MEMORY_21__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__18_ (.CK(CTS_52),
	.D(n_547),
	.Q(DPATH_RF_MEMORY_21__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__19_ (.CK(CTS_26),
	.D(n_546),
	.Q(DPATH_RF_MEMORY_21__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__20_ (.CK(CTS_21),
	.D(n_544),
	.Q(DPATH_RF_MEMORY_21__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__21_ (.CK(CTS_42),
	.D(n_542),
	.Q(DPATH_RF_MEMORY_21__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__22_ (.CK(CTS_42),
	.D(n_540),
	.Q(DPATH_RF_MEMORY_21__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__23_ (.CK(CTS_21),
	.D(n_538),
	.Q(DPATH_RF_MEMORY_21__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__24_ (.CK(CTS_51),
	.D(n_537),
	.Q(DPATH_RF_MEMORY_21__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__25_ (.CK(CTS_28),
	.D(n_536),
	.Q(DPATH_RF_MEMORY_21__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__26_ (.CK(CTS_9),
	.D(n_534),
	.Q(DPATH_RF_MEMORY_21__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__27_ (.CK(CTS_13),
	.D(n_533),
	.Q(DPATH_RF_MEMORY_21__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__28_ (.CK(CTS_29),
	.D(n_531),
	.Q(DPATH_RF_MEMORY_21__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__29_ (.CK(CTS_52),
	.D(n_529),
	.Q(DPATH_RF_MEMORY_21__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__30_ (.CK(CTS_51),
	.D(n_528),
	.Q(DPATH_RF_MEMORY_21__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_21__31_ (.CK(CTS_17),
	.D(n_526),
	.Q(DPATH_RF_MEMORY_21__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__0_ (.CK(CTS_18),
	.D(n_1146),
	.Q(DPATH_RF_MEMORY_22__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__1_ (.CK(CTS_16),
	.D(n_1145),
	.Q(DPATH_RF_MEMORY_22__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__2_ (.CK(CTS_50),
	.D(n_185),
	.Q(DPATH_RF_MEMORY_22__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__3_ (.CK(CTS_22),
	.D(n_1144),
	.Q(DPATH_RF_MEMORY_22__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__4_ (.CK(CTS_29),
	.D(n_1143),
	.Q(DPATH_RF_MEMORY_22__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__5_ (.CK(CTS_16),
	.D(n_1142),
	.Q(DPATH_RF_MEMORY_22__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__6_ (.CK(CTS_15),
	.D(n_1141),
	.Q(DPATH_RF_MEMORY_22__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__7_ (.CK(CTS_1),
	.D(n_1140),
	.Q(DPATH_RF_MEMORY_22__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__8_ (.CK(CTS_18),
	.D(n_1139),
	.Q(DPATH_RF_MEMORY_22__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__9_ (.CK(CTS_15),
	.D(n_1138),
	.Q(DPATH_RF_MEMORY_22__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__10_ (.CK(CTS_50),
	.D(n_1137),
	.Q(DPATH_RF_MEMORY_22__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__11_ (.CK(CTS_52),
	.D(n_1136),
	.Q(DPATH_RF_MEMORY_22__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__12_ (.CK(CTS_9),
	.D(n_1135),
	.Q(DPATH_RF_MEMORY_22__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__13_ (.CK(CTS_41),
	.D(n_1134),
	.Q(DPATH_RF_MEMORY_22__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__14_ (.CK(CTS_45),
	.D(n_1133),
	.Q(DPATH_RF_MEMORY_22__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__15_ (.CK(CTS_26),
	.D(n_1132),
	.Q(DPATH_RF_MEMORY_22__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__16_ (.CK(CTS_45),
	.D(n_1131),
	.Q(DPATH_RF_MEMORY_22__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__17_ (.CK(CTS_28),
	.D(n_1130),
	.Q(DPATH_RF_MEMORY_22__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__18_ (.CK(CTS_52),
	.D(n_1129),
	.Q(DPATH_RF_MEMORY_22__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__19_ (.CK(CTS_13),
	.D(n_1128),
	.Q(DPATH_RF_MEMORY_22__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__20_ (.CK(CTS_13),
	.D(n_1127),
	.Q(DPATH_RF_MEMORY_22__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__21_ (.CK(CTS_42),
	.D(n_1126),
	.Q(DPATH_RF_MEMORY_22__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__22_ (.CK(CTS_42),
	.D(n_1125),
	.Q(DPATH_RF_MEMORY_22__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__23_ (.CK(CTS_21),
	.D(n_1124),
	.Q(DPATH_RF_MEMORY_22__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__24_ (.CK(CTS_43),
	.D(n_1123),
	.Q(DPATH_RF_MEMORY_22__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__25_ (.CK(CTS_13),
	.D(n_1122),
	.Q(DPATH_RF_MEMORY_22__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__26_ (.CK(CTS_9),
	.D(n_1121),
	.Q(DPATH_RF_MEMORY_22__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__27_ (.CK(CTS_13),
	.D(n_1120),
	.Q(DPATH_RF_MEMORY_22__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__28_ (.CK(CTS_59),
	.D(n_1119),
	.Q(DPATH_RF_MEMORY_22__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__29_ (.CK(CTS_51),
	.D(n_1118),
	.Q(DPATH_RF_MEMORY_22__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__30_ (.CK(CTS_51),
	.D(n_1117),
	.Q(DPATH_RF_MEMORY_22__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_22__31_ (.CK(CTS_17),
	.D(n_1116),
	.Q(DPATH_RF_MEMORY_22__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__0_ (.CK(CTS_15),
	.D(n_464),
	.Q(DPATH_RF_MEMORY_23__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__1_ (.CK(CTS_16),
	.D(n_463),
	.Q(DPATH_RF_MEMORY_23__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__2_ (.CK(CTS_11),
	.D(n_163),
	.Q(DPATH_RF_MEMORY_23__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__3_ (.CK(CTS_1),
	.D(n_462),
	.Q(DPATH_RF_MEMORY_23__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__4_ (.CK(CTS_10),
	.D(n_461),
	.Q(DPATH_RF_MEMORY_23__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__5_ (.CK(CTS_14),
	.D(n_460),
	.Q(DPATH_RF_MEMORY_23__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__6_ (.CK(CTS_15),
	.D(n_459),
	.Q(DPATH_RF_MEMORY_23__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__7_ (.CK(CTS_1),
	.D(n_458),
	.Q(DPATH_RF_MEMORY_23__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__8_ (.CK(CTS_15),
	.D(n_457),
	.Q(DPATH_RF_MEMORY_23__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__9_ (.CK(CTS_1),
	.D(n_456),
	.Q(DPATH_RF_MEMORY_23__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__10_ (.CK(CTS_14),
	.D(n_455),
	.Q(DPATH_RF_MEMORY_23__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__11_ (.CK(CTS_52),
	.D(n_454),
	.Q(DPATH_RF_MEMORY_23__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__12_ (.CK(CTS_59),
	.D(n_453),
	.Q(DPATH_RF_MEMORY_23__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__13_ (.CK(CTS_14),
	.D(n_452),
	.Q(DPATH_RF_MEMORY_23__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__14_ (.CK(CTS_2),
	.D(n_451),
	.Q(DPATH_RF_MEMORY_23__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__15_ (.CK(CTS_37),
	.D(n_450),
	.Q(DPATH_RF_MEMORY_23__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__16_ (.CK(CTS_43),
	.D(n_449),
	.Q(DPATH_RF_MEMORY_23__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__17_ (.CK(CTS_38),
	.D(n_448),
	.Q(DPATH_RF_MEMORY_23__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__18_ (.CK(CTS_37),
	.D(n_447),
	.Q(DPATH_RF_MEMORY_23__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__19_ (.CK(CTS_35),
	.D(n_446),
	.Q(DPATH_RF_MEMORY_23__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__20_ (.CK(CTS_30),
	.D(n_445),
	.Q(DPATH_RF_MEMORY_23__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__21_ (.CK(CTS_52),
	.D(n_444),
	.Q(DPATH_RF_MEMORY_23__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__22_ (.CK(CTS_2),
	.D(n_443),
	.Q(DPATH_RF_MEMORY_23__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__23_ (.CK(CTS_34),
	.D(n_442),
	.Q(DPATH_RF_MEMORY_23__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__24_ (.CK(CTS_52),
	.D(n_441),
	.Q(DPATH_RF_MEMORY_23__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__25_ (.CK(CTS_26),
	.D(n_440),
	.Q(DPATH_RF_MEMORY_23__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__26_ (.CK(CTS_9),
	.D(n_439),
	.Q(DPATH_RF_MEMORY_23__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__27_ (.CK(CTS_34),
	.D(n_438),
	.Q(DPATH_RF_MEMORY_23__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__28_ (.CK(CTS_30),
	.D(n_437),
	.Q(DPATH_RF_MEMORY_23__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__29_ (.CK(CTS_51),
	.D(n_436),
	.Q(DPATH_RF_MEMORY_23__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__30_ (.CK(CTS_51),
	.D(n_435),
	.Q(DPATH_RF_MEMORY_23__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_23__31_ (.CK(CTS_33),
	.D(n_434),
	.Q(DPATH_RF_MEMORY_23__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__0_ (.CK(CTS_15),
	.D(n_1115),
	.Q(DPATH_RF_MEMORY_24__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__1_ (.CK(CTS_16),
	.D(n_1114),
	.Q(DPATH_RF_MEMORY_24__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__2_ (.CK(CTS_14),
	.D(n_184),
	.Q(DPATH_RF_MEMORY_24__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__3_ (.CK(CTS_1),
	.D(n_1113),
	.Q(DPATH_RF_MEMORY_24__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__4_ (.CK(CTS_33),
	.D(n_1112),
	.Q(DPATH_RF_MEMORY_24__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__5_ (.CK(CTS_14),
	.D(n_1111),
	.Q(DPATH_RF_MEMORY_24__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__6_ (.CK(CTS_4),
	.D(n_1110),
	.Q(DPATH_RF_MEMORY_24__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__7_ (.CK(CTS_5),
	.D(n_1109),
	.Q(DPATH_RF_MEMORY_24__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__8_ (.CK(CTS_15),
	.D(n_1108),
	.Q(DPATH_RF_MEMORY_24__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__9_ (.CK(CTS_1),
	.D(n_1107),
	.Q(DPATH_RF_MEMORY_24__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__10_ (.CK(CTS_14),
	.D(n_1106),
	.Q(DPATH_RF_MEMORY_24__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__11_ (.CK(CTS_52),
	.D(n_1105),
	.Q(DPATH_RF_MEMORY_24__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__12_ (.CK(CTS_9),
	.D(n_1104),
	.Q(DPATH_RF_MEMORY_24__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__13_ (.CK(CTS_14),
	.D(n_1103),
	.Q(DPATH_RF_MEMORY_24__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__14_ (.CK(CTS_2),
	.D(n_1102),
	.Q(DPATH_RF_MEMORY_24__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__15_ (.CK(CTS_35),
	.D(n_1101),
	.Q(DPATH_RF_MEMORY_24__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__16_ (.CK(CTS_42),
	.D(n_1100),
	.Q(DPATH_RF_MEMORY_24__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__17_ (.CK(CTS_26),
	.D(n_1099),
	.Q(DPATH_RF_MEMORY_24__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__18_ (.CK(CTS_35),
	.D(n_1098),
	.Q(DPATH_RF_MEMORY_24__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__19_ (.CK(CTS_34),
	.D(n_1097),
	.Q(DPATH_RF_MEMORY_24__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__20_ (.CK(CTS_30),
	.D(n_1096),
	.Q(DPATH_RF_MEMORY_24__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__21_ (.CK(CTS_51),
	.D(n_1095),
	.Q(DPATH_RF_MEMORY_24__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__22_ (.CK(CTS_2),
	.D(n_1094),
	.Q(DPATH_RF_MEMORY_24__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__23_ (.CK(CTS_34),
	.D(n_1093),
	.Q(DPATH_RF_MEMORY_24__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__24_ (.CK(CTS_52),
	.D(n_1092),
	.Q(DPATH_RF_MEMORY_24__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__25_ (.CK(CTS_35),
	.D(n_1091),
	.Q(DPATH_RF_MEMORY_24__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__26_ (.CK(CTS_9),
	.D(n_1090),
	.Q(DPATH_RF_MEMORY_24__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__27_ (.CK(CTS_34),
	.D(n_1089),
	.Q(DPATH_RF_MEMORY_24__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__28_ (.CK(CTS_30),
	.D(n_1088),
	.Q(DPATH_RF_MEMORY_24__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__29_ (.CK(CTS_44),
	.D(n_1087),
	.Q(DPATH_RF_MEMORY_24__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__30_ (.CK(CTS_51),
	.D(n_1086),
	.Q(DPATH_RF_MEMORY_24__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_24__31_ (.CK(CTS_33),
	.D(n_1085),
	.Q(DPATH_RF_MEMORY_24__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__0_ (.CK(CTS_4),
	.D(n_1084),
	.Q(DPATH_RF_MEMORY_25__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__1_ (.CK(CTS_17),
	.D(n_1083),
	.Q(DPATH_RF_MEMORY_25__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__2_ (.CK(CTS_10),
	.D(n_183),
	.Q(DPATH_RF_MEMORY_25__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__3_ (.CK(CTS_5),
	.D(n_1082),
	.Q(DPATH_RF_MEMORY_25__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__4_ (.CK(CTS_33),
	.D(n_1081),
	.Q(DPATH_RF_MEMORY_25__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__5_ (.CK(CTS_10),
	.D(n_1080),
	.Q(DPATH_RF_MEMORY_25__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__6_ (.CK(CTS_4),
	.D(n_1079),
	.Q(DPATH_RF_MEMORY_25__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__7_ (.CK(CTS_3),
	.D(n_1078),
	.Q(DPATH_RF_MEMORY_25__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__8_ (.CK(CTS_59),
	.D(n_1077),
	.Q(DPATH_RF_MEMORY_25__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__9_ (.CK(CTS_3),
	.D(n_1076),
	.Q(DPATH_RF_MEMORY_25__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__10_ (.CK(CTS_10),
	.D(n_1075),
	.Q(DPATH_RF_MEMORY_25__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__11_ (.CK(CTS_30),
	.D(n_1074),
	.Q(DPATH_RF_MEMORY_25__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__12_ (.CK(CTS_59),
	.D(n_1073),
	.Q(DPATH_RF_MEMORY_25__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__13_ (.CK(CTS_33),
	.D(n_1072),
	.Q(DPATH_RF_MEMORY_25__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__14_ (.CK(CTS_2),
	.D(n_1071),
	.Q(DPATH_RF_MEMORY_25__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__15_ (.CK(CTS_35),
	.D(n_1070),
	.Q(DPATH_RF_MEMORY_25__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__16_ (.CK(CTS_43),
	.D(n_1069),
	.Q(DPATH_RF_MEMORY_25__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__17_ (.CK(CTS_8),
	.D(n_1068),
	.Q(DPATH_RF_MEMORY_25__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__18_ (.CK(CTS_36),
	.D(n_1067),
	.Q(DPATH_RF_MEMORY_25__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__19_ (.CK(CTS_35),
	.D(n_1066),
	.Q(DPATH_RF_MEMORY_25__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__20_ (.CK(CTS_13),
	.D(n_1065),
	.Q(DPATH_RF_MEMORY_25__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__21_ (.CK(CTS_44),
	.D(n_1064),
	.Q(DPATH_RF_MEMORY_25__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__22_ (.CK(CTS_43),
	.D(n_1063),
	.Q(DPATH_RF_MEMORY_25__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__23_ (.CK(CTS_34),
	.D(n_1062),
	.Q(DPATH_RF_MEMORY_25__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__24_ (.CK(CTS_30),
	.D(n_1061),
	.Q(DPATH_RF_MEMORY_25__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__25_ (.CK(CTS_36),
	.D(n_1060),
	.Q(DPATH_RF_MEMORY_25__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__26_ (.CK(CTS_9),
	.D(n_1059),
	.Q(DPATH_RF_MEMORY_25__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__27_ (.CK(CTS_34),
	.D(n_1058),
	.Q(DPATH_RF_MEMORY_25__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__28_ (.CK(CTS_29),
	.D(n_1056),
	.Q(DPATH_RF_MEMORY_25__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__29_ (.CK(CTS_44),
	.D(n_1055),
	.Q(DPATH_RF_MEMORY_25__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__30_ (.CK(CTS_44),
	.D(n_1054),
	.Q(DPATH_RF_MEMORY_25__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_25__31_ (.CK(CTS_33),
	.D(n_1053),
	.Q(DPATH_RF_MEMORY_25__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__0_ (.CK(CTS_4),
	.D(n_1052),
	.Q(DPATH_RF_MEMORY_26__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__1_ (.CK(CTS_17),
	.D(n_1051),
	.Q(DPATH_RF_MEMORY_26__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__2_ (.CK(CTS_10),
	.D(n_182),
	.Q(DPATH_RF_MEMORY_26__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__3_ (.CK(CTS_5),
	.D(n_1050),
	.Q(DPATH_RF_MEMORY_26__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__4_ (.CK(CTS_33),
	.D(n_1049),
	.Q(DPATH_RF_MEMORY_26__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__5_ (.CK(CTS_10),
	.D(n_1048),
	.Q(DPATH_RF_MEMORY_26__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__6_ (.CK(CTS_4),
	.D(n_1047),
	.Q(DPATH_RF_MEMORY_26__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__7_ (.CK(CTS_3),
	.D(n_1046),
	.Q(DPATH_RF_MEMORY_26__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__8_ (.CK(CTS_3),
	.D(n_1045),
	.Q(DPATH_RF_MEMORY_26__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__9_ (.CK(CTS_3),
	.D(n_1044),
	.Q(DPATH_RF_MEMORY_26__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__10_ (.CK(CTS_10),
	.D(n_1043),
	.Q(DPATH_RF_MEMORY_26__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__11_ (.CK(CTS_30),
	.D(n_1042),
	.Q(DPATH_RF_MEMORY_26__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__12_ (.CK(CTS_59),
	.D(n_1041),
	.Q(DPATH_RF_MEMORY_26__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__13_ (.CK(CTS_33),
	.D(n_1039),
	.Q(DPATH_RF_MEMORY_26__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__14_ (.CK(CTS_2),
	.D(n_1038),
	.Q(DPATH_RF_MEMORY_26__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__15_ (.CK(CTS_35),
	.D(n_1036),
	.Q(DPATH_RF_MEMORY_26__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__16_ (.CK(CTS_43),
	.D(n_1035),
	.Q(DPATH_RF_MEMORY_26__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__17_ (.CK(CTS_8),
	.D(n_1034),
	.Q(DPATH_RF_MEMORY_26__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__18_ (.CK(CTS_34),
	.D(n_1033),
	.Q(DPATH_RF_MEMORY_26__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__19_ (.CK(CTS_35),
	.D(n_1031),
	.Q(DPATH_RF_MEMORY_26__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__20_ (.CK(CTS_30),
	.D(n_1029),
	.Q(DPATH_RF_MEMORY_26__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__21_ (.CK(CTS_44),
	.D(n_1027),
	.Q(DPATH_RF_MEMORY_26__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__22_ (.CK(CTS_43),
	.D(n_1026),
	.Q(DPATH_RF_MEMORY_26__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__23_ (.CK(CTS_34),
	.D(n_1025),
	.Q(DPATH_RF_MEMORY_26__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__24_ (.CK(CTS_30),
	.D(n_1023),
	.Q(DPATH_RF_MEMORY_26__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__25_ (.CK(CTS_36),
	.D(n_1022),
	.Q(DPATH_RF_MEMORY_26__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__26_ (.CK(CTS_9),
	.D(n_1020),
	.Q(DPATH_RF_MEMORY_26__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__27_ (.CK(CTS_34),
	.D(n_1018),
	.Q(DPATH_RF_MEMORY_26__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__28_ (.CK(CTS_29),
	.D(n_1017),
	.Q(DPATH_RF_MEMORY_26__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__29_ (.CK(CTS_44),
	.D(n_1015),
	.Q(DPATH_RF_MEMORY_26__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__30_ (.CK(CTS_44),
	.D(n_1014),
	.Q(DPATH_RF_MEMORY_26__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_26__31_ (.CK(CTS_33),
	.D(n_1013),
	.Q(DPATH_RF_MEMORY_26__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__0_ (.CK(CTS_15),
	.D(n_650),
	.Q(DPATH_RF_MEMORY_27__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__1_ (.CK(CTS_16),
	.D(n_649),
	.Q(DPATH_RF_MEMORY_27__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__2_ (.CK(CTS_10),
	.D(n_169),
	.Q(DPATH_RF_MEMORY_27__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__3_ (.CK(CTS_1),
	.D(n_648),
	.Q(DPATH_RF_MEMORY_27__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__4_ (.CK(CTS_10),
	.D(n_647),
	.Q(DPATH_RF_MEMORY_27__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__5_ (.CK(CTS_14),
	.D(n_646),
	.Q(DPATH_RF_MEMORY_27__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__6_ (.CK(CTS_15),
	.D(n_645),
	.Q(DPATH_RF_MEMORY_27__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__7_ (.CK(CTS_1),
	.D(n_644),
	.Q(DPATH_RF_MEMORY_27__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__8_ (.CK(CTS_15),
	.D(n_643),
	.Q(DPATH_RF_MEMORY_27__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__9_ (.CK(CTS_1),
	.D(n_642),
	.Q(DPATH_RF_MEMORY_27__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__10_ (.CK(CTS_14),
	.D(n_641),
	.Q(DPATH_RF_MEMORY_27__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__11_ (.CK(CTS_52),
	.D(n_640),
	.Q(DPATH_RF_MEMORY_27__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__12_ (.CK(CTS_43),
	.D(n_639),
	.Q(DPATH_RF_MEMORY_27__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__13_ (.CK(CTS_14),
	.D(n_638),
	.Q(DPATH_RF_MEMORY_27__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__14_ (.CK(CTS_43),
	.D(n_637),
	.Q(DPATH_RF_MEMORY_27__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__15_ (.CK(CTS_35),
	.D(n_636),
	.Q(DPATH_RF_MEMORY_27__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__16_ (.CK(CTS_43),
	.D(n_635),
	.Q(DPATH_RF_MEMORY_27__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__17_ (.CK(CTS_26),
	.D(n_634),
	.Q(DPATH_RF_MEMORY_27__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__18_ (.CK(CTS_35),
	.D(n_633),
	.Q(DPATH_RF_MEMORY_27__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__19_ (.CK(CTS_35),
	.D(n_632),
	.Q(DPATH_RF_MEMORY_27__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__20_ (.CK(CTS_30),
	.D(n_631),
	.Q(DPATH_RF_MEMORY_27__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__21_ (.CK(CTS_51),
	.D(n_630),
	.Q(DPATH_RF_MEMORY_27__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__22_ (.CK(CTS_43),
	.D(n_629),
	.Q(DPATH_RF_MEMORY_27__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__23_ (.CK(CTS_33),
	.D(n_628),
	.Q(DPATH_RF_MEMORY_27__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__24_ (.CK(CTS_52),
	.D(n_627),
	.Q(DPATH_RF_MEMORY_27__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__25_ (.CK(CTS_26),
	.D(n_626),
	.Q(DPATH_RF_MEMORY_27__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__26_ (.CK(CTS_9),
	.D(n_625),
	.Q(DPATH_RF_MEMORY_27__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__27_ (.CK(CTS_34),
	.D(n_624),
	.Q(DPATH_RF_MEMORY_27__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__28_ (.CK(CTS_21),
	.D(n_623),
	.Q(DPATH_RF_MEMORY_27__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__29_ (.CK(CTS_51),
	.D(n_622),
	.Q(DPATH_RF_MEMORY_27__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__30_ (.CK(CTS_51),
	.D(n_621),
	.Q(DPATH_RF_MEMORY_27__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_27__31_ (.CK(CTS_33),
	.D(n_620),
	.Q(DPATH_RF_MEMORY_27__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__0_ (.CK(CTS_4),
	.D(n_994),
	.Q(DPATH_RF_MEMORY_28__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__1_ (.CK(CTS_16),
	.D(n_993),
	.Q(DPATH_RF_MEMORY_28__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__2_ (.CK(CTS_10),
	.D(n_180),
	.Q(DPATH_RF_MEMORY_28__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__3_ (.CK(CTS_1),
	.D(n_991),
	.Q(DPATH_RF_MEMORY_28__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__4_ (.CK(CTS_10),
	.D(n_703),
	.Q(DPATH_RF_MEMORY_28__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__5_ (.CK(CTS_10),
	.D(n_988),
	.Q(DPATH_RF_MEMORY_28__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__6_ (.CK(CTS_15),
	.D(n_987),
	.Q(DPATH_RF_MEMORY_28__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__7_ (.CK(CTS_1),
	.D(n_986),
	.Q(DPATH_RF_MEMORY_28__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__8_ (.CK(CTS_15),
	.D(n_723),
	.Q(DPATH_RF_MEMORY_28__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__9_ (.CK(CTS_3),
	.D(n_984),
	.Q(DPATH_RF_MEMORY_28__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__10_ (.CK(CTS_10),
	.D(n_983),
	.Q(DPATH_RF_MEMORY_28__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__11_ (.CK(CTS_13),
	.D(n_982),
	.Q(DPATH_RF_MEMORY_28__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__12_ (.CK(CTS_9),
	.D(n_981),
	.Q(DPATH_RF_MEMORY_28__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__13_ (.CK(CTS_10),
	.D(n_980),
	.Q(DPATH_RF_MEMORY_28__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__14_ (.CK(CTS_43),
	.D(n_978),
	.Q(DPATH_RF_MEMORY_28__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__15_ (.CK(CTS_35),
	.D(n_977),
	.Q(DPATH_RF_MEMORY_28__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__16_ (.CK(CTS_43),
	.D(n_976),
	.Q(DPATH_RF_MEMORY_28__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__17_ (.CK(CTS_26),
	.D(n_975),
	.Q(DPATH_RF_MEMORY_28__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__18_ (.CK(CTS_35),
	.D(n_974),
	.Q(DPATH_RF_MEMORY_28__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__19_ (.CK(CTS_34),
	.D(n_973),
	.Q(DPATH_RF_MEMORY_28__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__20_ (.CK(CTS_13),
	.D(n_972),
	.Q(DPATH_RF_MEMORY_28__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__21_ (.CK(CTS_51),
	.D(n_971),
	.Q(DPATH_RF_MEMORY_28__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__22_ (.CK(CTS_43),
	.D(n_970),
	.Q(DPATH_RF_MEMORY_28__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__23_ (.CK(CTS_34),
	.D(n_969),
	.Q(DPATH_RF_MEMORY_28__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__24_ (.CK(CTS_52),
	.D(n_968),
	.Q(DPATH_RF_MEMORY_28__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__25_ (.CK(CTS_26),
	.D(n_967),
	.Q(DPATH_RF_MEMORY_28__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__26_ (.CK(CTS_9),
	.D(n_966),
	.Q(DPATH_RF_MEMORY_28__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__27_ (.CK(CTS_36),
	.D(n_965),
	.Q(DPATH_RF_MEMORY_28__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__28_ (.CK(CTS_29),
	.D(n_964),
	.Q(DPATH_RF_MEMORY_28__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__29_ (.CK(CTS_51),
	.D(n_963),
	.Q(DPATH_RF_MEMORY_28__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__30_ (.CK(CTS_51),
	.D(n_962),
	.Q(DPATH_RF_MEMORY_28__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_28__31_ (.CK(CTS_33),
	.D(n_961),
	.Q(DPATH_RF_MEMORY_28__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__0_ (.CK(CTS_4),
	.D(n_960),
	.Q(DPATH_RF_MEMORY_29__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__1_ (.CK(CTS_4),
	.D(n_959),
	.Q(DPATH_RF_MEMORY_29__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__2_ (.CK(CTS_14),
	.D(n_179),
	.Q(DPATH_RF_MEMORY_29__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__3_ (.CK(CTS_5),
	.D(n_958),
	.Q(DPATH_RF_MEMORY_29__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__4_ (.CK(CTS_33),
	.D(n_957),
	.Q(DPATH_RF_MEMORY_29__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__5_ (.CK(CTS_14),
	.D(n_955),
	.Q(DPATH_RF_MEMORY_29__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__6_ (.CK(CTS_4),
	.D(n_954),
	.Q(DPATH_RF_MEMORY_29__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__7_ (.CK(CTS_5),
	.D(n_953),
	.Q(DPATH_RF_MEMORY_29__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__8_ (.CK(CTS_59),
	.D(n_952),
	.Q(DPATH_RF_MEMORY_29__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__9_ (.CK(CTS_3),
	.D(n_951),
	.Q(DPATH_RF_MEMORY_29__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__10_ (.CK(CTS_10),
	.D(n_950),
	.Q(DPATH_RF_MEMORY_29__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__11_ (.CK(CTS_13),
	.D(n_949),
	.Q(DPATH_RF_MEMORY_29__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__12_ (.CK(CTS_59),
	.D(n_948),
	.Q(DPATH_RF_MEMORY_29__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__13_ (.CK(CTS_33),
	.D(n_947),
	.Q(DPATH_RF_MEMORY_29__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__14_ (.CK(CTS_2),
	.D(n_946),
	.Q(DPATH_RF_MEMORY_29__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__15_ (.CK(CTS_35),
	.D(n_945),
	.Q(DPATH_RF_MEMORY_29__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__16_ (.CK(CTS_42),
	.D(n_944),
	.Q(DPATH_RF_MEMORY_29__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__17_ (.CK(CTS_8),
	.D(n_943),
	.Q(DPATH_RF_MEMORY_29__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__18_ (.CK(CTS_35),
	.D(n_942),
	.Q(DPATH_RF_MEMORY_29__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__19_ (.CK(CTS_34),
	.D(n_941),
	.Q(DPATH_RF_MEMORY_29__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__20_ (.CK(CTS_13),
	.D(n_940),
	.Q(DPATH_RF_MEMORY_29__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__21_ (.CK(CTS_44),
	.D(n_939),
	.Q(DPATH_RF_MEMORY_29__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__22_ (.CK(CTS_2),
	.D(n_938),
	.Q(DPATH_RF_MEMORY_29__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__23_ (.CK(CTS_33),
	.D(n_937),
	.Q(DPATH_RF_MEMORY_29__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__24_ (.CK(CTS_30),
	.D(n_936),
	.Q(DPATH_RF_MEMORY_29__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__25_ (.CK(CTS_35),
	.D(n_935),
	.Q(DPATH_RF_MEMORY_29__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__26_ (.CK(CTS_9),
	.D(n_934),
	.Q(DPATH_RF_MEMORY_29__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__27_ (.CK(CTS_34),
	.D(n_933),
	.Q(DPATH_RF_MEMORY_29__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__28_ (.CK(CTS_21),
	.D(n_932),
	.Q(DPATH_RF_MEMORY_29__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__29_ (.CK(CTS_44),
	.D(n_931),
	.Q(DPATH_RF_MEMORY_29__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__30_ (.CK(CTS_44),
	.D(n_930),
	.Q(DPATH_RF_MEMORY_29__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_29__31_ (.CK(CTS_33),
	.D(n_929),
	.Q(DPATH_RF_MEMORY_29__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__0_ (.CK(CTS_4),
	.D(n_928),
	.Q(DPATH_RF_MEMORY_30__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__1_ (.CK(CTS_4),
	.D(n_927),
	.Q(DPATH_RF_MEMORY_30__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__2_ (.CK(CTS_14),
	.D(n_178),
	.Q(DPATH_RF_MEMORY_30__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__3_ (.CK(CTS_5),
	.D(n_926),
	.Q(DPATH_RF_MEMORY_30__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__4_ (.CK(CTS_33),
	.D(n_925),
	.Q(DPATH_RF_MEMORY_30__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__5_ (.CK(CTS_10),
	.D(n_924),
	.Q(DPATH_RF_MEMORY_30__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__6_ (.CK(CTS_4),
	.D(n_923),
	.Q(DPATH_RF_MEMORY_30__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__7_ (.CK(CTS_5),
	.D(n_922),
	.Q(DPATH_RF_MEMORY_30__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__8_ (.CK(CTS_4),
	.D(n_921),
	.Q(DPATH_RF_MEMORY_30__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__9_ (.CK(CTS_3),
	.D(n_920),
	.Q(DPATH_RF_MEMORY_30__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__10_ (.CK(CTS_10),
	.D(n_919),
	.Q(DPATH_RF_MEMORY_30__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__11_ (.CK(CTS_13),
	.D(n_918),
	.Q(DPATH_RF_MEMORY_30__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__12_ (.CK(CTS_59),
	.D(n_916),
	.Q(DPATH_RF_MEMORY_30__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__13_ (.CK(CTS_14),
	.D(n_915),
	.Q(DPATH_RF_MEMORY_30__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__14_ (.CK(CTS_2),
	.D(n_913),
	.Q(DPATH_RF_MEMORY_30__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__15_ (.CK(CTS_35),
	.D(n_912),
	.Q(DPATH_RF_MEMORY_30__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__16_ (.CK(CTS_42),
	.D(n_911),
	.Q(DPATH_RF_MEMORY_30__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__17_ (.CK(CTS_8),
	.D(n_910),
	.Q(DPATH_RF_MEMORY_30__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__18_ (.CK(CTS_35),
	.D(n_908),
	.Q(DPATH_RF_MEMORY_30__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__19_ (.CK(CTS_34),
	.D(n_956),
	.Q(DPATH_RF_MEMORY_30__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__20_ (.CK(CTS_13),
	.D(n_905),
	.Q(DPATH_RF_MEMORY_30__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__21_ (.CK(CTS_44),
	.D(n_904),
	.Q(DPATH_RF_MEMORY_30__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__22_ (.CK(CTS_2),
	.D(n_903),
	.Q(DPATH_RF_MEMORY_30__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__23_ (.CK(CTS_34),
	.D(n_996),
	.Q(DPATH_RF_MEMORY_30__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__24_ (.CK(CTS_30),
	.D(n_901),
	.Q(DPATH_RF_MEMORY_30__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__25_ (.CK(CTS_8),
	.D(n_899),
	.Q(DPATH_RF_MEMORY_30__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__26_ (.CK(CTS_9),
	.D(n_897),
	.Q(DPATH_RF_MEMORY_30__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__27_ (.CK(CTS_34),
	.D(n_896),
	.Q(DPATH_RF_MEMORY_30__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__28_ (.CK(CTS_30),
	.D(n_894),
	.Q(DPATH_RF_MEMORY_30__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__29_ (.CK(CTS_44),
	.D(n_893),
	.Q(DPATH_RF_MEMORY_30__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__30_ (.CK(CTS_44),
	.D(n_892),
	.Q(DPATH_RF_MEMORY_30__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_30__31_ (.CK(CTS_33),
	.D(n_1057),
	.Q(DPATH_RF_MEMORY_30__31_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__0_ (.CK(CTS_15),
	.D(n_619),
	.Q(DPATH_RF_MEMORY_31__0_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__1_ (.CK(CTS_16),
	.D(n_618),
	.Q(DPATH_RF_MEMORY_31__1_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__2_ (.CK(CTS_41),
	.D(n_168),
	.Q(DPATH_RF_MEMORY_31__2_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__3_ (.CK(CTS_22),
	.D(n_617),
	.Q(DPATH_RF_MEMORY_31__3_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__4_ (.CK(CTS_29),
	.D(n_616),
	.Q(DPATH_RF_MEMORY_31__4_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__5_ (.CK(CTS_16),
	.D(n_615),
	.Q(DPATH_RF_MEMORY_31__5_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__6_ (.CK(CTS_15),
	.D(n_614),
	.Q(DPATH_RF_MEMORY_31__6_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__7_ (.CK(CTS_22),
	.D(n_613),
	.Q(DPATH_RF_MEMORY_31__7_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__8_ (.CK(CTS_22),
	.D(n_612),
	.Q(DPATH_RF_MEMORY_31__8_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__9_ (.CK(CTS_1),
	.D(n_611),
	.Q(DPATH_RF_MEMORY_31__9_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__10_ (.CK(CTS_41),
	.D(n_610),
	.Q(DPATH_RF_MEMORY_31__10_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__11_ (.CK(CTS_52),
	.D(n_609),
	.Q(DPATH_RF_MEMORY_31__11_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__12_ (.CK(CTS_59),
	.D(n_608),
	.Q(DPATH_RF_MEMORY_31__12_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__13_ (.CK(CTS_40),
	.D(n_607),
	.Q(DPATH_RF_MEMORY_31__13_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__14_ (.CK(CTS_43),
	.D(n_606),
	.Q(DPATH_RF_MEMORY_31__14_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__15_ (.CK(CTS_26),
	.D(n_605),
	.Q(DPATH_RF_MEMORY_31__15_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__16_ (.CK(CTS_43),
	.D(n_604),
	.Q(DPATH_RF_MEMORY_31__16_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__17_ (.CK(CTS_28),
	.D(n_603),
	.Q(DPATH_RF_MEMORY_31__17_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__18_ (.CK(CTS_13),
	.D(n_602),
	.Q(DPATH_RF_MEMORY_31__18_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__19_ (.CK(CTS_26),
	.D(n_601),
	.Q(DPATH_RF_MEMORY_31__19_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__20_ (.CK(CTS_21),
	.D(n_600),
	.Q(DPATH_RF_MEMORY_31__20_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__21_ (.CK(CTS_43),
	.D(n_599),
	.Q(DPATH_RF_MEMORY_31__21_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__22_ (.CK(CTS_42),
	.D(n_598),
	.Q(DPATH_RF_MEMORY_31__22_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__23_ (.CK(CTS_8),
	.D(n_597),
	.Q(DPATH_RF_MEMORY_31__23_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__24_ (.CK(CTS_51),
	.D(n_596),
	.Q(DPATH_RF_MEMORY_31__24_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__25_ (.CK(CTS_13),
	.D(n_595),
	.Q(DPATH_RF_MEMORY_31__25_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__26_ (.CK(CTS_9),
	.D(n_594),
	.Q(DPATH_RF_MEMORY_31__26_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__27_ (.CK(CTS_8),
	.D(n_593),
	.Q(DPATH_RF_MEMORY_31__27_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__28_ (.CK(CTS_59),
	.D(n_592),
	.Q(DPATH_RF_MEMORY_31__28_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__29_ (.CK(CTS_51),
	.D(n_591),
	.Q(DPATH_RF_MEMORY_31__29_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__30_ (.CK(CTS_51),
	.D(n_590),
	.Q(DPATH_RF_MEMORY_31__30_));
   DFFQ_X2_50_SVT DPATH_RF_MEMORY_reg_31__31_ (.CK(CTS_32),
	.D(n_589),
	.Q(DPATH_RF_MEMORY_31__31_));
   NAND2_A_OAI21_X2_50_SVT g44075 (.A0N(DPATH_RF_MEMORY_22__0_),
	.A1N(n_72),
	.B0(FE_OFN93_n_117),
	.B1(n_72),
	.Q(n_1146));
   NAND2_A_OAI21_X2_50_SVT g44076 (.A0N(DPATH_RF_MEMORY_22__1_),
	.A1N(n_72),
	.B0(FE_OFN108_n_140),
	.B1(n_72),
	.Q(n_1145));
   NAND2_A_OAI21_X2_50_SVT g44077 (.A0N(DPATH_RF_MEMORY_22__3_),
	.A1N(n_72),
	.B0(FE_OFN111_n_144),
	.B1(n_72),
	.Q(n_1144));
   NAND2_A_OAI21_X2_50_SVT g44078 (.A0N(DPATH_RF_MEMORY_22__4_),
	.A1N(n_72),
	.B0(FE_OFN82_n_93),
	.B1(n_72),
	.Q(n_1143));
   NAND2_A_OAI21_X2_50_SVT g44079 (.A0N(DPATH_RF_MEMORY_22__5_),
	.A1N(n_72),
	.B0(FE_OFN116_n_152),
	.B1(n_72),
	.Q(n_1142));
   NAND2_A_OAI21_X2_50_SVT g44080 (.A0N(DPATH_RF_MEMORY_22__6_),
	.A1N(n_72),
	.B0(FE_OFN107_n_138),
	.B1(n_72),
	.Q(n_1141));
   NAND2_A_OAI21_X2_50_SVT g44081 (.A0N(DPATH_RF_MEMORY_22__7_),
	.A1N(n_72),
	.B0(FE_OFN88_n_107),
	.B1(n_72),
	.Q(n_1140));
   NAND2_A_OAI21_X2_50_SVT g44082 (.A0N(DPATH_RF_MEMORY_22__8_),
	.A1N(n_72),
	.B0(FE_OFN106_n_136),
	.B1(n_72),
	.Q(n_1139));
   NAND2_A_OAI21_X2_50_SVT g44083 (.A0N(DPATH_RF_MEMORY_22__9_),
	.A1N(n_72),
	.B0(FE_OFN96_n_121),
	.B1(n_72),
	.Q(n_1138));
   NAND2_A_OAI21_X2_50_SVT g44084 (.A0N(DPATH_RF_MEMORY_22__10_),
	.A1N(n_72),
	.B0(FE_OFN105_n_134),
	.B1(n_72),
	.Q(n_1137));
   NAND2_A_OAI21_X2_50_SVT g44085 (.A0N(DPATH_RF_MEMORY_22__11_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN74_n_72),
	.Q(n_1136));
   NAND2_A_OAI21_X2_50_SVT g44086 (.A0N(DPATH_RF_MEMORY_22__12_),
	.A1N(n_72),
	.B0(FE_OFN102_n_130),
	.B1(n_72),
	.Q(n_1135));
   NAND2_A_OAI21_X2_50_SVT g44087 (.A0N(DPATH_RF_MEMORY_22__13_),
	.A1N(n_72),
	.B0(FE_OFN110_n_142),
	.B1(n_72),
	.Q(n_1134));
   NAND2_A_OAI21_X2_50_SVT g44088 (.A0N(DPATH_RF_MEMORY_22__14_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN74_n_72),
	.Q(n_1133));
   NAND2_A_OAI21_X2_50_SVT g44089 (.A0N(DPATH_RF_MEMORY_22__15_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN74_n_72),
	.Q(n_1132));
   NAND2_A_OAI21_X2_50_SVT g44090 (.A0N(DPATH_RF_MEMORY_22__16_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN74_n_72),
	.Q(n_1131));
   NAND2_A_OAI21_X2_50_SVT g44091 (.A0N(DPATH_RF_MEMORY_22__17_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN74_n_72),
	.Q(n_1130));
   NAND2_A_OAI21_X2_50_SVT g44092 (.A0N(DPATH_RF_MEMORY_22__18_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN74_n_72),
	.Q(n_1129));
   NAND2_A_OAI21_X2_50_SVT g44093 (.A0N(DPATH_RF_MEMORY_22__19_),
	.A1N(n_72),
	.B0(FE_OFN92_n_115),
	.B1(n_72),
	.Q(n_1128));
   NAND2_A_OAI21_X2_50_SVT g44094 (.A0N(DPATH_RF_MEMORY_22__20_),
	.A1N(n_72),
	.B0(FE_OFN91_n_113),
	.B1(n_72),
	.Q(n_1127));
   NAND2_A_OAI21_X2_50_SVT g44095 (.A0N(DPATH_RF_MEMORY_22__21_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN74_n_72),
	.Q(n_1126));
   NAND2_A_OAI21_X2_50_SVT g44096 (.A0N(DPATH_RF_MEMORY_22__22_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN74_n_72),
	.Q(n_1125));
   NAND2_A_OAI21_X2_50_SVT g44097 (.A0N(DPATH_RF_MEMORY_22__23_),
	.A1N(n_72),
	.B0(FE_OFN97_n_123),
	.B1(n_72),
	.Q(n_1124));
   NAND2_A_OAI21_X2_50_SVT g44098 (.A0N(DPATH_RF_MEMORY_22__24_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN74_n_72),
	.Q(n_1123));
   NAND2_A_OAI21_X2_50_SVT g44099 (.A0N(DPATH_RF_MEMORY_22__25_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN74_n_72),
	.Q(n_1122));
   NAND2_A_OAI21_X2_50_SVT g44100 (.A0N(DPATH_RF_MEMORY_22__26_),
	.A1N(n_72),
	.B0(FE_OFN87_n_105),
	.B1(n_72),
	.Q(n_1121));
   NAND2_A_OAI21_X2_50_SVT g44101 (.A0N(DPATH_RF_MEMORY_22__27_),
	.A1N(n_72),
	.B0(FE_OFN86_n_103),
	.B1(n_72),
	.Q(n_1120));
   NAND2_A_OAI21_X2_50_SVT g44102 (.A0N(DPATH_RF_MEMORY_22__28_),
	.A1N(n_72),
	.B0(FE_OFN85_n_101),
	.B1(n_72),
	.Q(n_1119));
   NAND2_A_OAI21_X2_50_SVT g44103 (.A0N(DPATH_RF_MEMORY_22__29_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN74_n_72),
	.Q(n_1118));
   NAND2_A_OAI21_X2_50_SVT g44104 (.A0N(DPATH_RF_MEMORY_22__30_),
	.A1N(FE_OFN74_n_72),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN74_n_72),
	.Q(n_1117));
   NAND2_A_OAI21_X2_50_SVT g44105 (.A0N(DPATH_RF_MEMORY_22__31_),
	.A1N(n_72),
	.B0(FE_OFN119_n_95),
	.B1(n_72),
	.Q(n_1116));
   NAND2_A_OAI21_X2_50_SVT g44106 (.A0N(DPATH_RF_MEMORY_24__0_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN81_n_86),
	.Q(n_1115));
   NAND2_A_OAI21_X2_50_SVT g44107 (.A0N(DPATH_RF_MEMORY_24__1_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN81_n_86),
	.Q(n_1114));
   NAND2_A_OAI21_X2_50_SVT g44108 (.A0N(DPATH_RF_MEMORY_24__3_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN81_n_86),
	.Q(n_1113));
   NAND2_A_OAI21_X2_50_SVT g44109 (.A0N(DPATH_RF_MEMORY_24__4_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN81_n_86),
	.Q(n_1112));
   NAND2_A_OAI21_X2_50_SVT g44110 (.A0N(DPATH_RF_MEMORY_24__5_),
	.A1N(n_86),
	.B0(FE_OFN116_n_152),
	.B1(n_86),
	.Q(n_1111));
   NAND2_A_OAI21_X2_50_SVT g44111 (.A0N(DPATH_RF_MEMORY_24__6_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN81_n_86),
	.Q(n_1110));
   NAND2_A_OAI21_X2_50_SVT g44112 (.A0N(DPATH_RF_MEMORY_24__7_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN81_n_86),
	.Q(n_1109));
   NAND2_A_OAI21_X2_50_SVT g44113 (.A0N(DPATH_RF_MEMORY_24__8_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN81_n_86),
	.Q(n_1108));
   NAND2_A_OAI21_X2_50_SVT g44114 (.A0N(DPATH_RF_MEMORY_24__9_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN81_n_86),
	.Q(n_1107));
   NAND2_A_OAI21_X2_50_SVT g44115 (.A0N(DPATH_RF_MEMORY_24__10_),
	.A1N(n_86),
	.B0(FE_OFN105_n_134),
	.B1(n_86),
	.Q(n_1106));
   NAND2_A_OAI21_X2_50_SVT g44116 (.A0N(DPATH_RF_MEMORY_24__11_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN81_n_86),
	.Q(n_1105));
   NAND2_A_OAI21_X2_50_SVT g44117 (.A0N(DPATH_RF_MEMORY_24__12_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN81_n_86),
	.Q(n_1104));
   NAND2_A_OAI21_X2_50_SVT g44118 (.A0N(DPATH_RF_MEMORY_24__13_),
	.A1N(n_86),
	.B0(FE_OFN110_n_142),
	.B1(n_86),
	.Q(n_1103));
   NAND2_A_OAI21_X2_50_SVT g44119 (.A0N(DPATH_RF_MEMORY_24__14_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN81_n_86),
	.Q(n_1102));
   NAND2_A_OAI21_X2_50_SVT g44120 (.A0N(DPATH_RF_MEMORY_24__15_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN81_n_86),
	.Q(n_1101));
   NAND2_A_OAI21_X2_50_SVT g44121 (.A0N(DPATH_RF_MEMORY_24__16_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN81_n_86),
	.Q(n_1100));
   NAND2_A_OAI21_X2_50_SVT g44122 (.A0N(DPATH_RF_MEMORY_24__17_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN81_n_86),
	.Q(n_1099));
   NAND2_A_OAI21_X2_50_SVT g44123 (.A0N(DPATH_RF_MEMORY_24__18_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN81_n_86),
	.Q(n_1098));
   NAND2_A_OAI21_X2_50_SVT g44124 (.A0N(DPATH_RF_MEMORY_24__19_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN81_n_86),
	.Q(n_1097));
   NAND2_A_OAI21_X2_50_SVT g44125 (.A0N(DPATH_RF_MEMORY_24__20_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN81_n_86),
	.Q(n_1096));
   NAND2_A_OAI21_X2_50_SVT g44126 (.A0N(DPATH_RF_MEMORY_24__21_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN81_n_86),
	.Q(n_1095));
   NAND2_A_OAI21_X2_50_SVT g44127 (.A0N(DPATH_RF_MEMORY_24__22_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN81_n_86),
	.Q(n_1094));
   NAND2_A_OAI21_X2_50_SVT g44128 (.A0N(DPATH_RF_MEMORY_24__23_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN81_n_86),
	.Q(n_1093));
   NAND2_A_OAI21_X2_50_SVT g44129 (.A0N(DPATH_RF_MEMORY_24__24_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN81_n_86),
	.Q(n_1092));
   NAND2_A_OAI21_X2_50_SVT g44130 (.A0N(DPATH_RF_MEMORY_24__25_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN81_n_86),
	.Q(n_1091));
   NAND2_A_OAI21_X2_50_SVT g44131 (.A0N(DPATH_RF_MEMORY_24__26_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN81_n_86),
	.Q(n_1090));
   NAND2_A_OAI21_X2_50_SVT g44132 (.A0N(DPATH_RF_MEMORY_24__27_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN81_n_86),
	.Q(n_1089));
   NAND2_A_OAI21_X2_50_SVT g44133 (.A0N(DPATH_RF_MEMORY_24__28_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN81_n_86),
	.Q(n_1088));
   NAND2_A_OAI21_X2_50_SVT g44134 (.A0N(DPATH_RF_MEMORY_24__29_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN81_n_86),
	.Q(n_1087));
   NAND2_A_OAI21_X2_50_SVT g44135 (.A0N(DPATH_RF_MEMORY_24__30_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN81_n_86),
	.Q(n_1086));
   NAND2_A_OAI21_X2_50_SVT g44136 (.A0N(DPATH_RF_MEMORY_24__31_),
	.A1N(FE_OFN81_n_86),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN81_n_86),
	.Q(n_1085));
   NAND2_A_OAI21_X2_50_SVT g44137 (.A0N(DPATH_RF_MEMORY_25__0_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN0_n_2),
	.Q(n_1084));
   NAND2_A_OAI21_X2_50_SVT g44138 (.A0N(DPATH_RF_MEMORY_25__1_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN0_n_2),
	.Q(n_1083));
   NAND2_A_OAI21_X2_50_SVT g44139 (.A0N(DPATH_RF_MEMORY_25__3_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN0_n_2),
	.Q(n_1082));
   NAND2_A_OAI21_X2_50_SVT g44140 (.A0N(DPATH_RF_MEMORY_25__4_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN0_n_2),
	.Q(n_1081));
   NAND2_A_OAI21_X2_50_SVT g44141 (.A0N(DPATH_RF_MEMORY_25__5_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN0_n_2),
	.Q(n_1080));
   NAND2_A_OAI21_X2_50_SVT g44142 (.A0N(DPATH_RF_MEMORY_25__6_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN0_n_2),
	.Q(n_1079));
   NAND2_A_OAI21_X2_50_SVT g44143 (.A0N(DPATH_RF_MEMORY_25__7_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN0_n_2),
	.Q(n_1078));
   NAND2_A_OAI21_X2_50_SVT g44144 (.A0N(DPATH_RF_MEMORY_25__8_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN0_n_2),
	.Q(n_1077));
   NAND2_A_OAI21_X2_50_SVT g44145 (.A0N(DPATH_RF_MEMORY_25__9_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN0_n_2),
	.Q(n_1076));
   NAND2_A_OAI21_X2_50_SVT g44146 (.A0N(DPATH_RF_MEMORY_25__10_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN0_n_2),
	.Q(n_1075));
   NAND2_A_OAI21_X2_50_SVT g44147 (.A0N(DPATH_RF_MEMORY_25__11_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN0_n_2),
	.Q(n_1074));
   NAND2_A_OAI21_X2_50_SVT g44148 (.A0N(DPATH_RF_MEMORY_25__12_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN0_n_2),
	.Q(n_1073));
   NAND2_A_OAI21_X2_50_SVT g44149 (.A0N(DPATH_RF_MEMORY_25__13_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN0_n_2),
	.Q(n_1072));
   NAND2_A_OAI21_X2_50_SVT g44150 (.A0N(DPATH_RF_MEMORY_25__14_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN0_n_2),
	.Q(n_1071));
   NAND2_A_OAI21_X2_50_SVT g44151 (.A0N(DPATH_RF_MEMORY_25__15_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN0_n_2),
	.Q(n_1070));
   NAND2_A_OAI21_X2_50_SVT g44152 (.A0N(DPATH_RF_MEMORY_25__16_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN0_n_2),
	.Q(n_1069));
   NAND2_A_OAI21_X2_50_SVT g44153 (.A0N(DPATH_RF_MEMORY_25__17_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN0_n_2),
	.Q(n_1068));
   NAND2_A_OAI21_X2_50_SVT g44154 (.A0N(DPATH_RF_MEMORY_25__18_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN0_n_2),
	.Q(n_1067));
   NAND2_A_OAI21_X2_50_SVT g44155 (.A0N(DPATH_RF_MEMORY_25__19_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN0_n_2),
	.Q(n_1066));
   NAND2_A_OAI21_X2_50_SVT g44156 (.A0N(DPATH_RF_MEMORY_25__20_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN0_n_2),
	.Q(n_1065));
   NAND2_A_OAI21_X2_50_SVT g44157 (.A0N(DPATH_RF_MEMORY_25__21_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN0_n_2),
	.Q(n_1064));
   NAND2_A_OAI21_X2_50_SVT g44158 (.A0N(DPATH_RF_MEMORY_25__22_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN0_n_2),
	.Q(n_1063));
   NAND2_A_OAI21_X2_50_SVT g44159 (.A0N(DPATH_RF_MEMORY_25__23_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN0_n_2),
	.Q(n_1062));
   NAND2_A_OAI21_X2_50_SVT g44160 (.A0N(DPATH_RF_MEMORY_25__24_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN0_n_2),
	.Q(n_1061));
   NAND2_A_OAI21_X2_50_SVT g44161 (.A0N(DPATH_RF_MEMORY_25__25_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN0_n_2),
	.Q(n_1060));
   NAND2_A_OAI21_X2_50_SVT g44162 (.A0N(DPATH_RF_MEMORY_25__26_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN0_n_2),
	.Q(n_1059));
   NAND2_A_OAI21_X2_50_SVT g44163 (.A0N(DPATH_RF_MEMORY_25__27_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN0_n_2),
	.Q(n_1058));
   NAND2_A_OAI21_X2_50_SVT g44164 (.A0N(DPATH_RF_MEMORY_30__31_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN78_n_79),
	.Q(n_1057));
   NAND2_A_OAI21_X2_50_SVT g44165 (.A0N(DPATH_RF_MEMORY_25__28_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN0_n_2),
	.Q(n_1056));
   NAND2_A_OAI21_X2_50_SVT g44166 (.A0N(DPATH_RF_MEMORY_25__29_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN0_n_2),
	.Q(n_1055));
   NAND2_A_OAI21_X2_50_SVT g44167 (.A0N(DPATH_RF_MEMORY_25__30_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN0_n_2),
	.Q(n_1054));
   NAND2_A_OAI21_X2_50_SVT g44168 (.A0N(DPATH_RF_MEMORY_25__31_),
	.A1N(FE_OFN0_n_2),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN0_n_2),
	.Q(n_1053));
   NAND2_A_OAI21_X2_50_SVT g44169 (.A0N(DPATH_RF_MEMORY_26__0_),
	.A1N(n_82),
	.B0(FE_OFN93_n_117),
	.B1(n_82),
	.Q(n_1052));
   NAND2_A_OAI21_X2_50_SVT g44170 (.A0N(DPATH_RF_MEMORY_26__1_),
	.A1N(n_82),
	.B0(FE_OFN108_n_140),
	.B1(n_82),
	.Q(n_1051));
   NAND2_A_OAI21_X2_50_SVT g44171 (.A0N(DPATH_RF_MEMORY_26__3_),
	.A1N(n_82),
	.B0(FE_OFN111_n_144),
	.B1(n_82),
	.Q(n_1050));
   NAND2_A_OAI21_X2_50_SVT g44172 (.A0N(DPATH_RF_MEMORY_26__4_),
	.A1N(n_82),
	.B0(FE_OFN82_n_93),
	.B1(n_82),
	.Q(n_1049));
   NAND2_A_OAI21_X2_50_SVT g44173 (.A0N(DPATH_RF_MEMORY_26__5_),
	.A1N(n_82),
	.B0(FE_OFN116_n_152),
	.B1(n_82),
	.Q(n_1048));
   NAND2_A_OAI21_X2_50_SVT g44174 (.A0N(DPATH_RF_MEMORY_26__6_),
	.A1N(n_82),
	.B0(FE_OFN107_n_138),
	.B1(n_82),
	.Q(n_1047));
   NAND2_A_OAI21_X2_50_SVT g44175 (.A0N(DPATH_RF_MEMORY_26__7_),
	.A1N(n_82),
	.B0(FE_OFN88_n_107),
	.B1(n_82),
	.Q(n_1046));
   NAND2_A_OAI21_X2_50_SVT g44176 (.A0N(DPATH_RF_MEMORY_26__8_),
	.A1N(n_82),
	.B0(FE_OFN106_n_136),
	.B1(n_82),
	.Q(n_1045));
   NAND2_A_OAI21_X2_50_SVT g44177 (.A0N(DPATH_RF_MEMORY_26__9_),
	.A1N(n_82),
	.B0(FE_OFN96_n_121),
	.B1(n_82),
	.Q(n_1044));
   NAND2_A_OAI21_X2_50_SVT g44178 (.A0N(DPATH_RF_MEMORY_26__10_),
	.A1N(n_82),
	.B0(FE_OFN105_n_134),
	.B1(n_82),
	.Q(n_1043));
   NAND2_A_OAI21_X2_50_SVT g44179 (.A0N(DPATH_RF_MEMORY_26__11_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN79_n_82),
	.Q(n_1042));
   NAND2_A_OAI21_X2_50_SVT g44180 (.A0N(DPATH_RF_MEMORY_26__12_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN102_n_130),
	.B1(n_82),
	.Q(n_1041));
   NAND2_A_OAI21_X2_50_SVT g44181 (.A0N(DPATH_RF_MEMORY_8__1_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN15_n_83),
	.Q(n_1040));
   NAND2_A_OAI21_X2_50_SVT g44182 (.A0N(DPATH_RF_MEMORY_26__13_),
	.A1N(n_82),
	.B0(FE_OFN110_n_142),
	.B1(n_82),
	.Q(n_1039));
   NAND2_A_OAI21_X2_50_SVT g44183 (.A0N(DPATH_RF_MEMORY_26__14_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN79_n_82),
	.Q(n_1038));
   NAND2_A_OAI21_X2_50_SVT g44184 (.A0N(DPATH_RF_MEMORY_8__0_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN15_n_83),
	.Q(n_1037));
   NAND2_A_OAI21_X2_50_SVT g44185 (.A0N(DPATH_RF_MEMORY_26__15_),
	.A1N(n_82),
	.B0(FE_OFN99_n_125),
	.B1(n_82),
	.Q(n_1036));
   NAND2_A_OAI21_X2_50_SVT g44186 (.A0N(DPATH_RF_MEMORY_26__16_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN79_n_82),
	.Q(n_1035));
   NAND2_A_OAI21_X2_50_SVT g44187 (.A0N(DPATH_RF_MEMORY_26__17_),
	.A1N(n_82),
	.B0(FE_OFN95_n_119),
	.B1(n_82),
	.Q(n_1034));
   NAND2_A_OAI21_X2_50_SVT g44188 (.A0N(DPATH_RF_MEMORY_26__18_),
	.A1N(n_82),
	.B0(FE_OFN113_n_148),
	.B1(n_82),
	.Q(n_1033));
   NAND2_A_OAI21_X2_50_SVT g44189 (.A0N(DPATH_RF_MEMORY_8__3_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN15_n_83),
	.Q(n_1032));
   NAND2_A_OAI21_X2_50_SVT g44190 (.A0N(DPATH_RF_MEMORY_26__19_),
	.A1N(n_82),
	.B0(FE_OFN92_n_115),
	.B1(n_82),
	.Q(n_1031));
   NAND2_A_OAI21_X2_50_SVT g44191 (.A0N(DPATH_RF_MEMORY_8__4_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN15_n_83),
	.Q(n_1030));
   NAND2_A_OAI21_X2_50_SVT g44192 (.A0N(DPATH_RF_MEMORY_26__20_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN79_n_82),
	.Q(n_1029));
   NAND2_A_OAI21_X2_50_SVT g44193 (.A0N(DPATH_RF_MEMORY_8__5_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN15_n_83),
	.Q(n_1028));
   NAND2_A_OAI21_X2_50_SVT g44194 (.A0N(DPATH_RF_MEMORY_26__21_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN79_n_82),
	.Q(n_1027));
   NAND2_A_OAI21_X2_50_SVT g44195 (.A0N(DPATH_RF_MEMORY_26__22_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN79_n_82),
	.Q(n_1026));
   NAND2_A_OAI21_X2_50_SVT g44196 (.A0N(DPATH_RF_MEMORY_26__23_),
	.A1N(n_82),
	.B0(FE_OFN97_n_123),
	.B1(n_82),
	.Q(n_1025));
   NAND2_A_OAI21_X2_50_SVT g44197 (.A0N(DPATH_RF_MEMORY_8__6_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN15_n_83),
	.Q(n_1024));
   NAND2_A_OAI21_X2_50_SVT g44198 (.A0N(DPATH_RF_MEMORY_26__24_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN79_n_82),
	.Q(n_1023));
   NAND2_A_OAI21_X2_50_SVT g44199 (.A0N(DPATH_RF_MEMORY_26__25_),
	.A1N(n_82),
	.B0(FE_OFN89_n_109),
	.B1(n_82),
	.Q(n_1022));
   NAND2_A_OAI21_X2_50_SVT g44200 (.A0N(DPATH_RF_MEMORY_8__7_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN15_n_83),
	.Q(n_1021));
   NAND2_A_OAI21_X2_50_SVT g44201 (.A0N(DPATH_RF_MEMORY_26__26_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN79_n_82),
	.Q(n_1020));
   NAND2_A_OAI21_X2_50_SVT g44202 (.A0N(DPATH_RF_MEMORY_8__8_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN15_n_83),
	.Q(n_1019));
   NAND2_A_OAI21_X2_50_SVT g44203 (.A0N(DPATH_RF_MEMORY_26__27_),
	.A1N(n_82),
	.B0(FE_OFN86_n_103),
	.B1(n_82),
	.Q(n_1018));
   NAND2_A_OAI21_X2_50_SVT g44204 (.A0N(DPATH_RF_MEMORY_26__28_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN79_n_82),
	.Q(n_1017));
   NAND2_A_OAI21_X2_50_SVT g44205 (.A0N(DPATH_RF_MEMORY_8__9_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN15_n_83),
	.Q(n_1016));
   NAND2_A_OAI21_X2_50_SVT g44206 (.A0N(DPATH_RF_MEMORY_26__29_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN79_n_82),
	.Q(n_1015));
   NAND2_A_OAI21_X2_50_SVT g44207 (.A0N(DPATH_RF_MEMORY_26__30_),
	.A1N(FE_OFN79_n_82),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN79_n_82),
	.Q(n_1014));
   NAND2_A_OAI21_X2_50_SVT g44208 (.A0N(DPATH_RF_MEMORY_26__31_),
	.A1N(n_82),
	.B0(FE_OFN119_n_95),
	.B1(n_82),
	.Q(n_1013));
   NAND2_A_OAI21_X2_50_SVT g44209 (.A0N(DPATH_RF_MEMORY_8__10_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN15_n_83),
	.Q(n_1012));
   NAND2_A_OAI21_X2_50_SVT g44210 (.A0N(DPATH_RF_MEMORY_8__11_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN15_n_83),
	.Q(n_1011));
   NAND2_A_OAI21_X2_50_SVT g44211 (.A0N(DPATH_RF_MEMORY_8__12_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN15_n_83),
	.Q(n_1010));
   NAND2_A_OAI21_X2_50_SVT g44212 (.A0N(DPATH_RF_MEMORY_8__13_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN15_n_83),
	.Q(n_1009));
   NAND2_A_OAI21_X2_50_SVT g44213 (.A0N(DPATH_RF_MEMORY_8__14_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN15_n_83),
	.Q(n_1008));
   NAND2_A_OAI21_X2_50_SVT g44214 (.A0N(DPATH_RF_MEMORY_8__17_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN15_n_83),
	.Q(n_1007));
   NAND2_A_OAI21_X2_50_SVT g44215 (.A0N(DPATH_RF_MEMORY_8__15_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN15_n_83),
	.Q(n_1006));
   NAND2_A_OAI21_X2_50_SVT g44216 (.A0N(DPATH_RF_MEMORY_8__16_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN15_n_83),
	.Q(n_1005));
   NAND2_A_OAI21_X2_50_SVT g44217 (.A0N(DPATH_RF_MEMORY_8__18_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN15_n_83),
	.Q(n_1004));
   NAND2_A_OAI21_X2_50_SVT g44218 (.A0N(DPATH_RF_MEMORY_8__19_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN15_n_83),
	.Q(n_1003));
   NAND2_A_OAI21_X2_50_SVT g44219 (.A0N(DPATH_RF_MEMORY_8__20_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN15_n_83),
	.Q(n_1002));
   NAND2_A_OAI21_X2_50_SVT g44220 (.A0N(DPATH_RF_MEMORY_8__21_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN15_n_83),
	.Q(n_1001));
   NAND2_A_OAI21_X2_50_SVT g44221 (.A0N(DPATH_RF_MEMORY_8__22_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN15_n_83),
	.Q(n_1000));
   NAND2_A_OAI21_X2_50_SVT g44222 (.A0N(DPATH_RF_MEMORY_8__23_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN15_n_83),
	.Q(n_999));
   NAND2_A_OAI21_X2_50_SVT g44223 (.A0N(DPATH_RF_MEMORY_8__24_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN15_n_83),
	.Q(n_998));
   NAND2_A_OAI21_X2_50_SVT g44224 (.A0N(DPATH_RF_MEMORY_8__25_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN15_n_83),
	.Q(n_997));
   NAND2_A_OAI21_X2_50_SVT g44225 (.A0N(DPATH_RF_MEMORY_30__23_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN78_n_79),
	.Q(n_996));
   NAND2_A_OAI21_X2_50_SVT g44226 (.A0N(DPATH_RF_MEMORY_8__26_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN15_n_83),
	.Q(n_995));
   NAND2_A_OAI21_X2_50_SVT g44227 (.A0N(DPATH_RF_MEMORY_28__0_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN80_n_85),
	.Q(n_994));
   NAND2_A_OAI21_X2_50_SVT g44228 (.A0N(DPATH_RF_MEMORY_28__1_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN80_n_85),
	.Q(n_993));
   NAND2_A_OAI21_X2_50_SVT g44229 (.A0N(DPATH_RF_MEMORY_8__27_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN15_n_83),
	.Q(n_992));
   NAND2_A_OAI21_X2_50_SVT g44230 (.A0N(DPATH_RF_MEMORY_28__3_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN80_n_85),
	.Q(n_991));
   NAND2_A_OAI21_X2_50_SVT g44231 (.A0N(DPATH_RF_MEMORY_8__28_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN15_n_83),
	.Q(n_990));
   NAND2_A_OAI21_X2_50_SVT g44232 (.A0N(DPATH_RF_MEMORY_8__29_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN15_n_83),
	.Q(n_989));
   NAND2_A_OAI21_X2_50_SVT g44233 (.A0N(DPATH_RF_MEMORY_28__5_),
	.A1N(n_85),
	.B0(FE_OFN116_n_152),
	.B1(n_85),
	.Q(n_988));
   NAND2_A_OAI21_X2_50_SVT g44234 (.A0N(DPATH_RF_MEMORY_28__6_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN80_n_85),
	.Q(n_987));
   NAND2_A_OAI21_X2_50_SVT g44235 (.A0N(DPATH_RF_MEMORY_28__7_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN80_n_85),
	.Q(n_986));
   NAND2_A_OAI21_X2_50_SVT g44236 (.A0N(DPATH_RF_MEMORY_8__30_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN15_n_83),
	.Q(n_985));
   NAND2_A_OAI21_X2_50_SVT g44237 (.A0N(DPATH_RF_MEMORY_28__9_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN80_n_85),
	.Q(n_984));
   NAND2_A_OAI21_X2_50_SVT g44238 (.A0N(DPATH_RF_MEMORY_28__10_),
	.A1N(n_85),
	.B0(FE_OFN105_n_134),
	.B1(n_85),
	.Q(n_983));
   NAND2_A_OAI21_X2_50_SVT g44239 (.A0N(DPATH_RF_MEMORY_28__11_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN80_n_85),
	.Q(n_982));
   NAND2_A_OAI21_X2_50_SVT g44240 (.A0N(DPATH_RF_MEMORY_28__12_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN80_n_85),
	.Q(n_981));
   NAND2_A_OAI21_X2_50_SVT g44241 (.A0N(DPATH_RF_MEMORY_28__13_),
	.A1N(n_85),
	.B0(FE_OFN110_n_142),
	.B1(n_85),
	.Q(n_980));
   NAND2_A_OAI21_X2_50_SVT g44242 (.A0N(DPATH_RF_MEMORY_8__31_),
	.A1N(FE_OFN15_n_83),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN15_n_83),
	.Q(n_979));
   NAND2_A_OAI21_X2_50_SVT g44243 (.A0N(DPATH_RF_MEMORY_28__14_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN80_n_85),
	.Q(n_978));
   NAND2_A_OAI21_X2_50_SVT g44244 (.A0N(DPATH_RF_MEMORY_28__15_),
	.A1N(n_85),
	.B0(FE_OFN99_n_125),
	.B1(n_85),
	.Q(n_977));
   NAND2_A_OAI21_X2_50_SVT g44245 (.A0N(DPATH_RF_MEMORY_28__16_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN80_n_85),
	.Q(n_976));
   NAND2_A_OAI21_X2_50_SVT g44246 (.A0N(DPATH_RF_MEMORY_28__17_),
	.A1N(n_85),
	.B0(FE_OFN95_n_119),
	.B1(n_85),
	.Q(n_975));
   NAND2_A_OAI21_X2_50_SVT g44247 (.A0N(DPATH_RF_MEMORY_28__18_),
	.A1N(n_85),
	.B0(FE_OFN113_n_148),
	.B1(n_85),
	.Q(n_974));
   NAND2_A_OAI21_X2_50_SVT g44248 (.A0N(DPATH_RF_MEMORY_28__19_),
	.A1N(n_85),
	.B0(FE_OFN92_n_115),
	.B1(n_85),
	.Q(n_973));
   NAND2_A_OAI21_X2_50_SVT g44249 (.A0N(DPATH_RF_MEMORY_28__20_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN80_n_85),
	.Q(n_972));
   NAND2_A_OAI21_X2_50_SVT g44250 (.A0N(DPATH_RF_MEMORY_28__21_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN80_n_85),
	.Q(n_971));
   NAND2_A_OAI21_X2_50_SVT g44251 (.A0N(DPATH_RF_MEMORY_28__22_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN80_n_85),
	.Q(n_970));
   NAND2_A_OAI21_X2_50_SVT g44252 (.A0N(DPATH_RF_MEMORY_28__23_),
	.A1N(n_85),
	.B0(FE_OFN97_n_123),
	.B1(n_85),
	.Q(n_969));
   NAND2_A_OAI21_X2_50_SVT g44253 (.A0N(DPATH_RF_MEMORY_28__24_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN80_n_85),
	.Q(n_968));
   NAND2_A_OAI21_X2_50_SVT g44254 (.A0N(DPATH_RF_MEMORY_28__25_),
	.A1N(n_85),
	.B0(FE_OFN89_n_109),
	.B1(n_85),
	.Q(n_967));
   NAND2_A_OAI21_X2_50_SVT g44255 (.A0N(DPATH_RF_MEMORY_28__26_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN80_n_85),
	.Q(n_966));
   NAND2_A_OAI21_X2_50_SVT g44256 (.A0N(DPATH_RF_MEMORY_28__27_),
	.A1N(n_85),
	.B0(FE_OFN86_n_103),
	.B1(n_85),
	.Q(n_965));
   NAND2_A_OAI21_X2_50_SVT g44257 (.A0N(DPATH_RF_MEMORY_28__28_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN80_n_85),
	.Q(n_964));
   NAND2_A_OAI21_X2_50_SVT g44258 (.A0N(DPATH_RF_MEMORY_28__29_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN80_n_85),
	.Q(n_963));
   NAND2_A_OAI21_X2_50_SVT g44259 (.A0N(DPATH_RF_MEMORY_28__30_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN80_n_85),
	.Q(n_962));
   NAND2_A_OAI21_X2_50_SVT g44260 (.A0N(DPATH_RF_MEMORY_28__31_),
	.A1N(n_85),
	.B0(FE_OFN119_n_95),
	.B1(n_85),
	.Q(n_961));
   NAND2_A_OAI21_X2_50_SVT g44261 (.A0N(DPATH_RF_MEMORY_29__0_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN4_n_67),
	.Q(n_960));
   NAND2_A_OAI21_X2_50_SVT g44262 (.A0N(DPATH_RF_MEMORY_29__1_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN4_n_67),
	.Q(n_959));
   NAND2_A_OAI21_X2_50_SVT g44263 (.A0N(DPATH_RF_MEMORY_29__3_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN4_n_67),
	.Q(n_958));
   NAND2_A_OAI21_X2_50_SVT g44264 (.A0N(DPATH_RF_MEMORY_29__4_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN4_n_67),
	.Q(n_957));
   NAND2_A_OAI21_X2_50_SVT g44265 (.A0N(DPATH_RF_MEMORY_30__19_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN78_n_79),
	.Q(n_956));
   NAND2_A_OAI21_X2_50_SVT g44266 (.A0N(DPATH_RF_MEMORY_29__5_),
	.A1N(n_67),
	.B0(FE_OFN116_n_152),
	.B1(n_67),
	.Q(n_955));
   NAND2_A_OAI21_X2_50_SVT g44267 (.A0N(DPATH_RF_MEMORY_29__6_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN4_n_67),
	.Q(n_954));
   NAND2_A_OAI21_X2_50_SVT g44268 (.A0N(DPATH_RF_MEMORY_29__7_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN4_n_67),
	.Q(n_953));
   NAND2_A_OAI21_X2_50_SVT g44269 (.A0N(DPATH_RF_MEMORY_29__8_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN4_n_67),
	.Q(n_952));
   NAND2_A_OAI21_X2_50_SVT g44270 (.A0N(DPATH_RF_MEMORY_29__9_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN4_n_67),
	.Q(n_951));
   NAND2_A_OAI21_X2_50_SVT g44271 (.A0N(DPATH_RF_MEMORY_29__10_),
	.A1N(n_67),
	.B0(FE_OFN105_n_134),
	.B1(n_67),
	.Q(n_950));
   NAND2_A_OAI21_X2_50_SVT g44272 (.A0N(DPATH_RF_MEMORY_29__11_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN4_n_67),
	.Q(n_949));
   NAND2_A_OAI21_X2_50_SVT g44273 (.A0N(DPATH_RF_MEMORY_29__12_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN4_n_67),
	.Q(n_948));
   NAND2_A_OAI21_X2_50_SVT g44274 (.A0N(DPATH_RF_MEMORY_29__13_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN4_n_67),
	.Q(n_947));
   NAND2_A_OAI21_X2_50_SVT g44275 (.A0N(DPATH_RF_MEMORY_29__14_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN4_n_67),
	.Q(n_946));
   NAND2_A_OAI21_X2_50_SVT g44276 (.A0N(DPATH_RF_MEMORY_29__15_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN4_n_67),
	.Q(n_945));
   NAND2_A_OAI21_X2_50_SVT g44277 (.A0N(DPATH_RF_MEMORY_29__16_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN4_n_67),
	.Q(n_944));
   NAND2_A_OAI21_X2_50_SVT g44278 (.A0N(DPATH_RF_MEMORY_29__17_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN4_n_67),
	.Q(n_943));
   NAND2_A_OAI21_X2_50_SVT g44279 (.A0N(DPATH_RF_MEMORY_29__18_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN4_n_67),
	.Q(n_942));
   NAND2_A_OAI21_X2_50_SVT g44280 (.A0N(DPATH_RF_MEMORY_29__19_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN4_n_67),
	.Q(n_941));
   NAND2_A_OAI21_X2_50_SVT g44281 (.A0N(DPATH_RF_MEMORY_29__20_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN4_n_67),
	.Q(n_940));
   NAND2_A_OAI21_X2_50_SVT g44282 (.A0N(DPATH_RF_MEMORY_29__21_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN4_n_67),
	.Q(n_939));
   NAND2_A_OAI21_X2_50_SVT g44283 (.A0N(DPATH_RF_MEMORY_29__22_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN4_n_67),
	.Q(n_938));
   NAND2_A_OAI21_X2_50_SVT g44284 (.A0N(DPATH_RF_MEMORY_29__23_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN4_n_67),
	.Q(n_937));
   NAND2_A_OAI21_X2_50_SVT g44285 (.A0N(DPATH_RF_MEMORY_29__24_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN4_n_67),
	.Q(n_936));
   NAND2_A_OAI21_X2_50_SVT g44286 (.A0N(DPATH_RF_MEMORY_29__25_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN4_n_67),
	.Q(n_935));
   NAND2_A_OAI21_X2_50_SVT g44287 (.A0N(DPATH_RF_MEMORY_29__26_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN4_n_67),
	.Q(n_934));
   NAND2_A_OAI21_X2_50_SVT g44288 (.A0N(DPATH_RF_MEMORY_29__27_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN4_n_67),
	.Q(n_933));
   NAND2_A_OAI21_X2_50_SVT g44289 (.A0N(DPATH_RF_MEMORY_29__28_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN4_n_67),
	.Q(n_932));
   NAND2_A_OAI21_X2_50_SVT g44290 (.A0N(DPATH_RF_MEMORY_29__29_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN4_n_67),
	.Q(n_931));
   NAND2_A_OAI21_X2_50_SVT g44291 (.A0N(DPATH_RF_MEMORY_29__30_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN4_n_67),
	.Q(n_930));
   NAND2_A_OAI21_X2_50_SVT g44292 (.A0N(DPATH_RF_MEMORY_29__31_),
	.A1N(FE_OFN4_n_67),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN4_n_67),
	.Q(n_929));
   NAND2_A_OAI21_X2_50_SVT g44293 (.A0N(DPATH_RF_MEMORY_30__0_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN78_n_79),
	.Q(n_928));
   NAND2_A_OAI21_X2_50_SVT g44294 (.A0N(DPATH_RF_MEMORY_30__1_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN78_n_79),
	.Q(n_927));
   NAND2_A_OAI21_X2_50_SVT g44295 (.A0N(DPATH_RF_MEMORY_30__3_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN78_n_79),
	.Q(n_926));
   NAND2_A_OAI21_X2_50_SVT g44296 (.A0N(DPATH_RF_MEMORY_30__4_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN78_n_79),
	.Q(n_925));
   NAND2_A_OAI21_X2_50_SVT g44297 (.A0N(DPATH_RF_MEMORY_30__5_),
	.A1N(n_79),
	.B0(FE_OFN116_n_152),
	.B1(n_79),
	.Q(n_924));
   NAND2_A_OAI21_X2_50_SVT g44298 (.A0N(DPATH_RF_MEMORY_30__6_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN78_n_79),
	.Q(n_923));
   NAND2_A_OAI21_X2_50_SVT g44299 (.A0N(DPATH_RF_MEMORY_30__7_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN78_n_79),
	.Q(n_922));
   NAND2_A_OAI21_X2_50_SVT g44300 (.A0N(DPATH_RF_MEMORY_30__8_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN78_n_79),
	.Q(n_921));
   NAND2_A_OAI21_X2_50_SVT g44301 (.A0N(DPATH_RF_MEMORY_30__9_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN78_n_79),
	.Q(n_920));
   NAND2_A_OAI21_X2_50_SVT g44302 (.A0N(DPATH_RF_MEMORY_30__10_),
	.A1N(n_79),
	.B0(FE_OFN105_n_134),
	.B1(n_79),
	.Q(n_919));
   NAND2_A_OAI21_X2_50_SVT g44303 (.A0N(DPATH_RF_MEMORY_30__11_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN78_n_79),
	.Q(n_918));
   NAND2_A_OAI21_X2_50_SVT g44304 (.A0N(DPATH_RF_MEMORY_10__1_),
	.A1N(n_81),
	.B0(FE_OFN108_n_140),
	.B1(n_81),
	.Q(n_917));
   NAND2_A_OAI21_X2_50_SVT g44305 (.A0N(DPATH_RF_MEMORY_30__12_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN78_n_79),
	.Q(n_916));
   NAND2_A_OAI21_X2_50_SVT g44306 (.A0N(DPATH_RF_MEMORY_30__13_),
	.A1N(n_79),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN78_n_79),
	.Q(n_915));
   NAND2_A_OAI21_X2_50_SVT g44307 (.A0N(DPATH_RF_MEMORY_10__0_),
	.A1N(n_81),
	.B0(FE_OFN93_n_117),
	.B1(n_81),
	.Q(n_914));
   NAND2_A_OAI21_X2_50_SVT g44308 (.A0N(DPATH_RF_MEMORY_30__14_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN78_n_79),
	.Q(n_913));
   NAND2_A_OAI21_X2_50_SVT g44309 (.A0N(DPATH_RF_MEMORY_30__15_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN78_n_79),
	.Q(n_912));
   NAND2_A_OAI21_X2_50_SVT g44310 (.A0N(DPATH_RF_MEMORY_30__16_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN78_n_79),
	.Q(n_911));
   NAND2_A_OAI21_X2_50_SVT g44311 (.A0N(DPATH_RF_MEMORY_30__17_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN78_n_79),
	.Q(n_910));
   NAND2_A_OAI21_X2_50_SVT g44312 (.A0N(DPATH_RF_MEMORY_10__3_),
	.A1N(n_81),
	.B0(FE_OFN111_n_144),
	.B1(n_81),
	.Q(n_909));
   NAND2_A_OAI21_X2_50_SVT g44313 (.A0N(DPATH_RF_MEMORY_30__18_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN78_n_79),
	.Q(n_908));
   NAND2_A_OAI21_X2_50_SVT g44314 (.A0N(DPATH_RF_MEMORY_10__4_),
	.A1N(n_81),
	.B0(FE_OFN82_n_93),
	.B1(n_81),
	.Q(n_907));
   NAND2_A_OAI21_X2_50_SVT g44315 (.A0N(DPATH_RF_MEMORY_10__5_),
	.A1N(n_81),
	.B0(FE_OFN116_n_152),
	.B1(n_81),
	.Q(n_906));
   NAND2_A_OAI21_X2_50_SVT g44316 (.A0N(DPATH_RF_MEMORY_30__20_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN78_n_79),
	.Q(n_905));
   NAND2_A_OAI21_X2_50_SVT g44317 (.A0N(DPATH_RF_MEMORY_30__21_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN78_n_79),
	.Q(n_904));
   NAND2_A_OAI21_X2_50_SVT g44318 (.A0N(DPATH_RF_MEMORY_30__22_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN78_n_79),
	.Q(n_903));
   NAND2_A_OAI21_X2_50_SVT g44319 (.A0N(DPATH_RF_MEMORY_10__6_),
	.A1N(n_81),
	.B0(FE_OFN107_n_138),
	.B1(n_81),
	.Q(n_902));
   NAND2_A_OAI21_X2_50_SVT g44320 (.A0N(DPATH_RF_MEMORY_30__24_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN78_n_79),
	.Q(n_901));
   NAND2_A_OAI21_X2_50_SVT g44321 (.A0N(DPATH_RF_MEMORY_10__7_),
	.A1N(n_81),
	.B0(FE_OFN88_n_107),
	.B1(n_81),
	.Q(n_900));
   NAND2_A_OAI21_X2_50_SVT g44322 (.A0N(DPATH_RF_MEMORY_30__25_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN78_n_79),
	.Q(n_899));
   NAND2_A_OAI21_X2_50_SVT g44323 (.A0N(DPATH_RF_MEMORY_10__8_),
	.A1N(n_81),
	.B0(FE_OFN106_n_136),
	.B1(n_81),
	.Q(n_898));
   NAND2_A_OAI21_X2_50_SVT g44324 (.A0N(DPATH_RF_MEMORY_30__26_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN78_n_79),
	.Q(n_897));
   NAND2_A_OAI21_X2_50_SVT g44325 (.A0N(DPATH_RF_MEMORY_30__27_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN78_n_79),
	.Q(n_896));
   NAND2_A_OAI21_X2_50_SVT g44326 (.A0N(DPATH_RF_MEMORY_10__9_),
	.A1N(n_81),
	.B0(FE_OFN96_n_121),
	.B1(n_81),
	.Q(n_895));
   NAND2_A_OAI21_X2_50_SVT g44327 (.A0N(DPATH_RF_MEMORY_30__28_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN78_n_79),
	.Q(n_894));
   NAND2_A_OAI21_X2_50_SVT g44328 (.A0N(DPATH_RF_MEMORY_30__29_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN78_n_79),
	.Q(n_893));
   NAND2_A_OAI21_X2_50_SVT g44329 (.A0N(DPATH_RF_MEMORY_30__30_),
	.A1N(FE_OFN78_n_79),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN78_n_79),
	.Q(n_892));
   NAND2_A_OAI21_X2_50_SVT g44330 (.A0N(DPATH_RF_MEMORY_10__10_),
	.A1N(n_81),
	.B0(FE_OFN105_n_134),
	.B1(n_81),
	.Q(n_891));
   NAND2_A_OAI21_X2_50_SVT g44331 (.A0N(DPATH_RF_MEMORY_10__11_),
	.A1N(n_81),
	.B0(FE_OFN103_n_132),
	.B1(n_81),
	.Q(n_890));
   NAND2_A_OAI21_X2_50_SVT g44332 (.A0N(DPATH_RF_MEMORY_10__12_),
	.A1N(n_81),
	.B0(FE_OFN102_n_130),
	.B1(n_81),
	.Q(n_889));
   NAND2_A_OAI21_X2_50_SVT g44333 (.A0N(DPATH_RF_MEMORY_10__13_),
	.A1N(n_81),
	.B0(FE_OFN110_n_142),
	.B1(n_81),
	.Q(n_888));
   NAND2_A_OAI21_X2_50_SVT g44334 (.A0N(DPATH_RF_MEMORY_10__14_),
	.A1N(n_81),
	.B0(FE_OFN100_n_127),
	.B1(n_81),
	.Q(n_887));
   NAND2_A_OAI21_X2_50_SVT g44335 (.A0N(DPATH_RF_MEMORY_10__15_),
	.A1N(n_81),
	.B0(FE_OFN99_n_125),
	.B1(n_81),
	.Q(n_886));
   NAND2_A_OAI21_X2_50_SVT g44336 (.A0N(DPATH_RF_MEMORY_10__16_),
	.A1N(n_81),
	.B0(FE_OFN117_n_154),
	.B1(n_81),
	.Q(n_885));
   NAND2_A_OAI21_X2_50_SVT g44337 (.A0N(DPATH_RF_MEMORY_10__17_),
	.A1N(n_81),
	.B0(FE_OFN95_n_119),
	.B1(n_81),
	.Q(n_884));
   NAND2_A_OAI21_X2_50_SVT g44338 (.A0N(DPATH_RF_MEMORY_10__18_),
	.A1N(n_81),
	.B0(FE_OFN113_n_148),
	.B1(n_81),
	.Q(n_883));
   NAND2_A_OAI21_X2_50_SVT g44339 (.A0N(DPATH_RF_MEMORY_10__19_),
	.A1N(n_81),
	.B0(FE_OFN92_n_115),
	.B1(n_81),
	.Q(n_882));
   NAND2_A_OAI21_X2_50_SVT g44340 (.A0N(DPATH_RF_MEMORY_10__20_),
	.A1N(n_81),
	.B0(FE_OFN91_n_113),
	.B1(n_81),
	.Q(n_881));
   NAND2_A_OAI21_X2_50_SVT g44341 (.A0N(DPATH_RF_MEMORY_10__21_),
	.A1N(n_81),
	.B0(FE_OFN112_n_146),
	.B1(n_81),
	.Q(n_880));
   NAND2_A_OAI21_X2_50_SVT g44342 (.A0N(DPATH_RF_MEMORY_10__22_),
	.A1N(n_81),
	.B0(FE_OFN114_n_150),
	.B1(n_81),
	.Q(n_879));
   NAND2_A_OAI21_X2_50_SVT g44343 (.A0N(DPATH_RF_MEMORY_10__23_),
	.A1N(n_81),
	.B0(FE_OFN97_n_123),
	.B1(n_81),
	.Q(n_878));
   NAND2_A_OAI21_X2_50_SVT g44344 (.A0N(DPATH_RF_MEMORY_10__24_),
	.A1N(n_81),
	.B0(FE_OFN90_n_111),
	.B1(n_81),
	.Q(n_877));
   NAND2_A_OAI21_X2_50_SVT g44345 (.A0N(DPATH_RF_MEMORY_10__25_),
	.A1N(n_81),
	.B0(FE_OFN89_n_109),
	.B1(n_81),
	.Q(n_876));
   NAND2_A_OAI21_X2_50_SVT g44346 (.A0N(DPATH_RF_MEMORY_10__26_),
	.A1N(n_81),
	.B0(FE_OFN87_n_105),
	.B1(n_81),
	.Q(n_875));
   NAND2_A_OAI21_X2_50_SVT g44347 (.A0N(DPATH_RF_MEMORY_10__27_),
	.A1N(n_81),
	.B0(FE_OFN86_n_103),
	.B1(n_81),
	.Q(n_874));
   NAND2_A_OAI21_X2_50_SVT g44348 (.A0N(DPATH_RF_MEMORY_10__28_),
	.A1N(n_81),
	.B0(FE_OFN85_n_101),
	.B1(n_81),
	.Q(n_873));
   NAND2_A_OAI21_X2_50_SVT g44349 (.A0N(DPATH_RF_MEMORY_10__29_),
	.A1N(n_81),
	.B0(FE_OFN84_n_99),
	.B1(n_81),
	.Q(n_872));
   NAND2_A_OAI21_X2_50_SVT g44350 (.A0N(DPATH_RF_MEMORY_10__30_),
	.A1N(n_81),
	.B0(FE_OFN83_n_97),
	.B1(n_81),
	.Q(n_871));
   NAND2_A_OAI21_X2_50_SVT g44351 (.A0N(DPATH_RF_MEMORY_10__31_),
	.A1N(n_81),
	.B0(FE_OFN119_n_95),
	.B1(n_81),
	.Q(n_870));
   NAND2_A_OAI21_X2_50_SVT g44352 (.A0N(DPATH_RF_MEMORY_12__0_),
	.A1N(n_62),
	.B0(FE_OFN93_n_117),
	.B1(n_62),
	.Q(n_869));
   NAND2_A_OAI21_X2_50_SVT g44353 (.A0N(DPATH_RF_MEMORY_12__1_),
	.A1N(n_62),
	.B0(FE_OFN108_n_140),
	.B1(n_62),
	.Q(n_868));
   NAND2_A_OAI21_X2_50_SVT g44354 (.A0N(DPATH_RF_MEMORY_12__3_),
	.A1N(n_62),
	.B0(FE_OFN111_n_144),
	.B1(n_62),
	.Q(n_867));
   NAND2_A_OAI21_X2_50_SVT g44355 (.A0N(DPATH_RF_MEMORY_12__4_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN82_n_93),
	.B1(n_62),
	.Q(n_866));
   NAND2_A_OAI21_X2_50_SVT g44356 (.A0N(DPATH_RF_MEMORY_12__5_),
	.A1N(n_62),
	.B0(FE_OFN116_n_152),
	.B1(n_62),
	.Q(n_865));
   NAND2_A_OAI21_X2_50_SVT g44357 (.A0N(DPATH_RF_MEMORY_12__6_),
	.A1N(n_62),
	.B0(FE_OFN107_n_138),
	.B1(n_62),
	.Q(n_864));
   NAND2_A_OAI21_X2_50_SVT g44358 (.A0N(DPATH_RF_MEMORY_12__7_),
	.A1N(n_62),
	.B0(FE_OFN88_n_107),
	.B1(n_62),
	.Q(n_863));
   NAND2_A_OAI21_X2_50_SVT g44359 (.A0N(DPATH_RF_MEMORY_12__8_),
	.A1N(n_62),
	.B0(FE_OFN106_n_136),
	.B1(n_62),
	.Q(n_862));
   NAND2_A_OAI21_X2_50_SVT g44360 (.A0N(DPATH_RF_MEMORY_12__9_),
	.A1N(n_62),
	.B0(FE_OFN96_n_121),
	.B1(n_62),
	.Q(n_861));
   NAND2_A_OAI21_X2_50_SVT g44361 (.A0N(DPATH_RF_MEMORY_12__10_),
	.A1N(n_62),
	.B0(FE_OFN105_n_134),
	.B1(n_62),
	.Q(n_860));
   NAND2_A_OAI21_X2_50_SVT g44362 (.A0N(DPATH_RF_MEMORY_12__11_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN2_n_62),
	.Q(n_859));
   NAND2_A_OAI21_X2_50_SVT g44363 (.A0N(DPATH_RF_MEMORY_12__12_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN2_n_62),
	.Q(n_858));
   NAND2_A_OAI21_X2_50_SVT g44364 (.A0N(DPATH_RF_MEMORY_12__13_),
	.A1N(n_62),
	.B0(FE_OFN110_n_142),
	.B1(n_62),
	.Q(n_857));
   NAND2_A_OAI21_X2_50_SVT g44365 (.A0N(DPATH_RF_MEMORY_12__14_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN2_n_62),
	.Q(n_856));
   NAND2_A_OAI21_X2_50_SVT g44366 (.A0N(DPATH_RF_MEMORY_12__15_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN2_n_62),
	.Q(n_855));
   NAND2_A_OAI21_X2_50_SVT g44367 (.A0N(DPATH_RF_MEMORY_12__16_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN2_n_62),
	.Q(n_854));
   NAND2_A_OAI21_X2_50_SVT g44368 (.A0N(DPATH_RF_MEMORY_12__17_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN2_n_62),
	.Q(n_853));
   NAND2_A_OAI21_X2_50_SVT g44369 (.A0N(DPATH_RF_MEMORY_12__18_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN2_n_62),
	.Q(n_852));
   NAND2_A_OAI21_X2_50_SVT g44370 (.A0N(DPATH_RF_MEMORY_12__19_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN2_n_62),
	.Q(n_851));
   NAND2_A_OAI21_X2_50_SVT g44371 (.A0N(DPATH_RF_MEMORY_12__20_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN2_n_62),
	.Q(n_850));
   NAND2_A_OAI21_X2_50_SVT g44372 (.A0N(DPATH_RF_MEMORY_12__21_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN2_n_62),
	.Q(n_849));
   NAND2_A_OAI21_X2_50_SVT g44373 (.A0N(DPATH_RF_MEMORY_12__22_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN2_n_62),
	.Q(n_848));
   NAND2_A_OAI21_X2_50_SVT g44374 (.A0N(DPATH_RF_MEMORY_12__23_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN2_n_62),
	.Q(n_847));
   NAND2_A_OAI21_X2_50_SVT g44375 (.A0N(DPATH_RF_MEMORY_12__24_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN2_n_62),
	.Q(n_846));
   NAND2_A_OAI21_X2_50_SVT g44376 (.A0N(DPATH_RF_MEMORY_12__25_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN2_n_62),
	.Q(n_845));
   NAND2_A_OAI21_X2_50_SVT g44377 (.A0N(DPATH_RF_MEMORY_12__26_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN2_n_62),
	.Q(n_844));
   NAND2_A_OAI21_X2_50_SVT g44378 (.A0N(DPATH_RF_MEMORY_12__27_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN2_n_62),
	.Q(n_843));
   NAND2_A_OAI21_X2_50_SVT g44379 (.A0N(DPATH_RF_MEMORY_12__28_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN2_n_62),
	.Q(n_842));
   NAND2_A_OAI21_X2_50_SVT g44380 (.A0N(DPATH_RF_MEMORY_12__29_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN2_n_62),
	.Q(n_841));
   NAND2_A_OAI21_X2_50_SVT g44381 (.A0N(DPATH_RF_MEMORY_12__30_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN2_n_62),
	.Q(n_840));
   NAND2_A_OAI21_X2_50_SVT g44382 (.A0N(DPATH_RF_MEMORY_12__31_),
	.A1N(FE_OFN2_n_62),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN2_n_62),
	.Q(n_839));
   NAND2_A_OAI21_X2_50_SVT g44383 (.A0N(DPATH_RF_MEMORY_14__0_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN5_n_69),
	.Q(n_838));
   NAND2_A_OAI21_X2_50_SVT g44384 (.A0N(DPATH_RF_MEMORY_14__1_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN5_n_69),
	.Q(n_837));
   NAND2_A_OAI21_X2_50_SVT g44385 (.A0N(DPATH_RF_MEMORY_14__3_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN5_n_69),
	.Q(n_836));
   NAND2_A_OAI21_X2_50_SVT g44386 (.A0N(DPATH_RF_MEMORY_14__4_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN5_n_69),
	.Q(n_835));
   NAND2_A_OAI21_X2_50_SVT g44387 (.A0N(DPATH_RF_MEMORY_14__5_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN5_n_69),
	.Q(n_834));
   NAND2_A_OAI21_X2_50_SVT g44388 (.A0N(DPATH_RF_MEMORY_14__6_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN5_n_69),
	.Q(n_833));
   NAND2_A_OAI21_X2_50_SVT g44389 (.A0N(DPATH_RF_MEMORY_14__7_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN5_n_69),
	.Q(n_832));
   NAND2_A_OAI21_X2_50_SVT g44390 (.A0N(DPATH_RF_MEMORY_14__8_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN5_n_69),
	.Q(n_831));
   NAND2_A_OAI21_X2_50_SVT g44391 (.A0N(DPATH_RF_MEMORY_14__9_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN5_n_69),
	.Q(n_830));
   NAND2_A_OAI21_X2_50_SVT g44392 (.A0N(DPATH_RF_MEMORY_14__10_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN5_n_69),
	.Q(n_829));
   NAND2_A_OAI21_X2_50_SVT g44393 (.A0N(DPATH_RF_MEMORY_14__11_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN5_n_69),
	.Q(n_828));
   NAND2_A_OAI21_X2_50_SVT g44394 (.A0N(DPATH_RF_MEMORY_14__12_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN5_n_69),
	.Q(n_827));
   NAND2_A_OAI21_X2_50_SVT g44395 (.A0N(DPATH_RF_MEMORY_14__13_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN5_n_69),
	.Q(n_826));
   NAND2_A_OAI21_X2_50_SVT g44396 (.A0N(DPATH_RF_MEMORY_14__14_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN5_n_69),
	.Q(n_825));
   NAND2_A_OAI21_X2_50_SVT g44397 (.A0N(DPATH_RF_MEMORY_14__15_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN5_n_69),
	.Q(n_824));
   NAND2_A_OAI21_X2_50_SVT g44398 (.A0N(DPATH_RF_MEMORY_14__16_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN5_n_69),
	.Q(n_823));
   NAND2_A_OAI21_X2_50_SVT g44399 (.A0N(DPATH_RF_MEMORY_14__17_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN5_n_69),
	.Q(n_822));
   NAND2_A_OAI21_X2_50_SVT g44400 (.A0N(DPATH_RF_MEMORY_14__18_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN5_n_69),
	.Q(n_821));
   NAND2_A_OAI21_X2_50_SVT g44401 (.A0N(DPATH_RF_MEMORY_14__19_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN5_n_69),
	.Q(n_820));
   NAND2_A_OAI21_X2_50_SVT g44402 (.A0N(DPATH_RF_MEMORY_14__20_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN5_n_69),
	.Q(n_819));
   NAND2_A_OAI21_X2_50_SVT g44403 (.A0N(DPATH_RF_MEMORY_14__21_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN5_n_69),
	.Q(n_818));
   NAND2_A_OAI21_X2_50_SVT g44404 (.A0N(DPATH_RF_MEMORY_14__22_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN5_n_69),
	.Q(n_817));
   NAND2_A_OAI21_X2_50_SVT g44405 (.A0N(DPATH_RF_MEMORY_14__23_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN5_n_69),
	.Q(n_816));
   NAND2_A_OAI21_X2_50_SVT g44406 (.A0N(DPATH_RF_MEMORY_14__24_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN5_n_69),
	.Q(n_815));
   NAND2_A_OAI21_X2_50_SVT g44407 (.A0N(DPATH_RF_MEMORY_14__25_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN5_n_69),
	.Q(n_814));
   NAND2_A_OAI21_X2_50_SVT g44408 (.A0N(DPATH_RF_MEMORY_14__26_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN5_n_69),
	.Q(n_813));
   NAND2_A_OAI21_X2_50_SVT g44409 (.A0N(DPATH_RF_MEMORY_14__27_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN5_n_69),
	.Q(n_812));
   NAND2_A_OAI21_X2_50_SVT g44410 (.A0N(DPATH_RF_MEMORY_14__28_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN5_n_69),
	.Q(n_811));
   NAND2_A_OAI21_X2_50_SVT g44411 (.A0N(DPATH_RF_MEMORY_14__29_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN5_n_69),
	.Q(n_810));
   NAND2_A_OAI21_X2_50_SVT g44412 (.A0N(DPATH_RF_MEMORY_14__30_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN5_n_69),
	.Q(n_809));
   NAND2_A_OAI21_X2_50_SVT g44413 (.A0N(DPATH_RF_MEMORY_14__31_),
	.A1N(FE_OFN5_n_69),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN5_n_69),
	.Q(n_808));
   NAND2_A_OAI21_X2_50_SVT g44414 (.A0N(DPATH_RF_MEMORY_16__0_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN75_n_73),
	.Q(n_807));
   NAND2_A_OAI21_X2_50_SVT g44415 (.A0N(DPATH_RF_MEMORY_16__1_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN75_n_73),
	.Q(n_806));
   NAND2_A_OAI21_X2_50_SVT g44416 (.A0N(DPATH_RF_MEMORY_16__3_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN75_n_73),
	.Q(n_805));
   NAND2_A_OAI21_X2_50_SVT g44417 (.A0N(DPATH_RF_MEMORY_16__4_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN75_n_73),
	.Q(n_804));
   NAND2_A_OAI21_X2_50_SVT g44418 (.A0N(DPATH_RF_MEMORY_16__5_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN75_n_73),
	.Q(n_803));
   NAND2_A_OAI21_X2_50_SVT g44419 (.A0N(DPATH_RF_MEMORY_16__6_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN75_n_73),
	.Q(n_802));
   NAND2_A_OAI21_X2_50_SVT g44420 (.A0N(DPATH_RF_MEMORY_16__7_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN75_n_73),
	.Q(n_801));
   NAND2_A_OAI21_X2_50_SVT g44421 (.A0N(DPATH_RF_MEMORY_16__8_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN75_n_73),
	.Q(n_800));
   NAND2_A_OAI21_X2_50_SVT g44422 (.A0N(DPATH_RF_MEMORY_16__9_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN75_n_73),
	.Q(n_799));
   NAND2_A_OAI21_X2_50_SVT g44423 (.A0N(DPATH_RF_MEMORY_16__10_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN75_n_73),
	.Q(n_798));
   NAND2_A_OAI21_X2_50_SVT g44424 (.A0N(DPATH_RF_MEMORY_16__11_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN75_n_73),
	.Q(n_797));
   NAND2_A_OAI21_X2_50_SVT g44425 (.A0N(DPATH_RF_MEMORY_16__12_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN75_n_73),
	.Q(n_796));
   NAND2_A_OAI21_X2_50_SVT g44426 (.A0N(DPATH_RF_MEMORY_16__13_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN75_n_73),
	.Q(n_795));
   NAND2_A_OAI21_X2_50_SVT g44427 (.A0N(DPATH_RF_MEMORY_16__14_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN75_n_73),
	.Q(n_794));
   NAND2_A_OAI21_X2_50_SVT g44428 (.A0N(DPATH_RF_MEMORY_16__15_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN75_n_73),
	.Q(n_793));
   NAND2_A_OAI21_X2_50_SVT g44429 (.A0N(DPATH_RF_MEMORY_16__16_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN75_n_73),
	.Q(n_792));
   NAND2_A_OAI21_X2_50_SVT g44430 (.A0N(DPATH_RF_MEMORY_16__17_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN75_n_73),
	.Q(n_791));
   NAND2_A_OAI21_X2_50_SVT g44431 (.A0N(DPATH_RF_MEMORY_16__18_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN75_n_73),
	.Q(n_790));
   NAND2_A_OAI21_X2_50_SVT g44432 (.A0N(DPATH_RF_MEMORY_16__19_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN75_n_73),
	.Q(n_789));
   NAND2_A_OAI21_X2_50_SVT g44433 (.A0N(DPATH_RF_MEMORY_16__20_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN75_n_73),
	.Q(n_788));
   NAND2_A_OAI21_X2_50_SVT g44434 (.A0N(DPATH_RF_MEMORY_16__21_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN75_n_73),
	.Q(n_787));
   NAND2_A_OAI21_X2_50_SVT g44435 (.A0N(DPATH_RF_MEMORY_16__22_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN75_n_73),
	.Q(n_786));
   NAND2_A_OAI21_X2_50_SVT g44436 (.A0N(DPATH_RF_MEMORY_16__23_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN75_n_73),
	.Q(n_785));
   NAND2_A_OAI21_X2_50_SVT g44437 (.A0N(DPATH_RF_MEMORY_16__24_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN75_n_73),
	.Q(n_784));
   NAND2_A_OAI21_X2_50_SVT g44438 (.A0N(DPATH_RF_MEMORY_16__25_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN75_n_73),
	.Q(n_783));
   NAND2_A_OAI21_X2_50_SVT g44439 (.A0N(DPATH_RF_MEMORY_16__26_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN75_n_73),
	.Q(n_782));
   NAND2_A_OAI21_X2_50_SVT g44440 (.A0N(DPATH_RF_MEMORY_16__27_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN75_n_73),
	.Q(n_781));
   NAND2_A_OAI21_X2_50_SVT g44441 (.A0N(DPATH_RF_MEMORY_16__28_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN75_n_73),
	.Q(n_780));
   NAND2_A_OAI21_X2_50_SVT g44442 (.A0N(DPATH_RF_MEMORY_16__29_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN75_n_73),
	.Q(n_779));
   NAND2_A_OAI21_X2_50_SVT g44443 (.A0N(DPATH_RF_MEMORY_16__30_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN75_n_73),
	.Q(n_778));
   NAND2_A_OAI21_X2_50_SVT g44444 (.A0N(DPATH_RF_MEMORY_16__31_),
	.A1N(FE_OFN75_n_73),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN75_n_73),
	.Q(n_777));
   NAND2_A_OAI21_X2_50_SVT g44445 (.A0N(DPATH_RF_MEMORY_18__0_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN76_n_75),
	.Q(n_776));
   NAND2_A_OAI21_X2_50_SVT g44446 (.A0N(DPATH_RF_MEMORY_18__1_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN76_n_75),
	.Q(n_775));
   NAND2_A_OAI21_X2_50_SVT g44447 (.A0N(DPATH_RF_MEMORY_18__3_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN76_n_75),
	.Q(n_774));
   NAND2_A_OAI21_X2_50_SVT g44448 (.A0N(DPATH_RF_MEMORY_18__4_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN76_n_75),
	.Q(n_773));
   NAND2_A_OAI21_X2_50_SVT g44449 (.A0N(DPATH_RF_MEMORY_18__5_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN76_n_75),
	.Q(n_772));
   NAND2_A_OAI21_X2_50_SVT g44450 (.A0N(DPATH_RF_MEMORY_18__6_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN76_n_75),
	.Q(n_771));
   NAND2_A_OAI21_X2_50_SVT g44451 (.A0N(DPATH_RF_MEMORY_18__7_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN76_n_75),
	.Q(n_770));
   NAND2_A_OAI21_X2_50_SVT g44452 (.A0N(DPATH_RF_MEMORY_4__0_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN3_n_64),
	.Q(n_769));
   NAND2_A_OAI21_X2_50_SVT g44453 (.A0N(DPATH_RF_MEMORY_18__8_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN76_n_75),
	.Q(n_768));
   NAND2_A_OAI21_X2_50_SVT g44454 (.A0N(DPATH_RF_MEMORY_18__9_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN76_n_75),
	.Q(n_767));
   NAND2_A_OAI21_X2_50_SVT g44455 (.A0N(DPATH_RF_MEMORY_18__10_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN76_n_75),
	.Q(n_766));
   NAND2_A_OAI21_X2_50_SVT g44456 (.A0N(DPATH_RF_MEMORY_18__11_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN76_n_75),
	.Q(n_765));
   NAND2_A_OAI21_X2_50_SVT g44457 (.A0N(DPATH_RF_MEMORY_18__12_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN76_n_75),
	.Q(n_764));
   NAND2_A_OAI21_X2_50_SVT g44458 (.A0N(DPATH_RF_MEMORY_18__13_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN76_n_75),
	.Q(n_763));
   NAND2_A_OAI21_X2_50_SVT g44459 (.A0N(DPATH_RF_MEMORY_18__14_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN76_n_75),
	.Q(n_762));
   NAND2_A_OAI21_X2_50_SVT g44460 (.A0N(DPATH_RF_MEMORY_18__15_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN76_n_75),
	.Q(n_761));
   NAND2_A_OAI21_X2_50_SVT g44461 (.A0N(DPATH_RF_MEMORY_4__3_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN3_n_64),
	.Q(n_760));
   NAND2_A_OAI21_X2_50_SVT g44462 (.A0N(DPATH_RF_MEMORY_18__16_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN76_n_75),
	.Q(n_759));
   NAND2_A_OAI21_X2_50_SVT g44463 (.A0N(DPATH_RF_MEMORY_18__17_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN76_n_75),
	.Q(n_758));
   NAND2_A_OAI21_X2_50_SVT g44464 (.A0N(DPATH_RF_MEMORY_4__1_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN108_n_140),
	.B1(FE_OFN3_n_64),
	.Q(n_757));
   NAND2_A_OAI21_X2_50_SVT g44465 (.A0N(DPATH_RF_MEMORY_4__4_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN3_n_64),
	.Q(n_756));
   NAND2_A_OAI21_X2_50_SVT g44466 (.A0N(DPATH_RF_MEMORY_18__18_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN76_n_75),
	.Q(n_755));
   NAND2_A_OAI21_X2_50_SVT g44467 (.A0N(DPATH_RF_MEMORY_18__19_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN76_n_75),
	.Q(n_754));
   NAND2_A_OAI21_X2_50_SVT g44468 (.A0N(DPATH_RF_MEMORY_18__20_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN76_n_75),
	.Q(n_753));
   NAND2_A_OAI21_X2_50_SVT g44469 (.A0N(DPATH_RF_MEMORY_18__21_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN76_n_75),
	.Q(n_752));
   NAND2_A_OAI21_X2_50_SVT g44470 (.A0N(DPATH_RF_MEMORY_4__5_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN116_n_152),
	.B1(FE_OFN3_n_64),
	.Q(n_751));
   NAND2_A_OAI21_X2_50_SVT g44471 (.A0N(DPATH_RF_MEMORY_4__6_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN107_n_138),
	.B1(FE_OFN3_n_64),
	.Q(n_750));
   NAND2_A_OAI21_X2_50_SVT g44472 (.A0N(DPATH_RF_MEMORY_18__22_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN76_n_75),
	.Q(n_749));
   NAND2_A_OAI21_X2_50_SVT g44473 (.A0N(DPATH_RF_MEMORY_18__23_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN76_n_75),
	.Q(n_748));
   NAND2_A_OAI21_X2_50_SVT g44474 (.A0N(DPATH_RF_MEMORY_4__7_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN3_n_64),
	.Q(n_747));
   NAND2_A_OAI21_X2_50_SVT g44475 (.A0N(DPATH_RF_MEMORY_18__24_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN76_n_75),
	.Q(n_746));
   NAND2_A_OAI21_X2_50_SVT g44476 (.A0N(DPATH_RF_MEMORY_18__25_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN76_n_75),
	.Q(n_745));
   NAND2_A_OAI21_X2_50_SVT g44477 (.A0N(DPATH_RF_MEMORY_4__8_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN3_n_64),
	.Q(n_744));
   NAND2_A_OAI21_X2_50_SVT g44478 (.A0N(DPATH_RF_MEMORY_18__26_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN76_n_75),
	.Q(n_743));
   NAND2_A_OAI21_X2_50_SVT g44479 (.A0N(DPATH_RF_MEMORY_18__27_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN76_n_75),
	.Q(n_742));
   NAND2_A_OAI21_X2_50_SVT g44480 (.A0N(DPATH_RF_MEMORY_18__28_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN76_n_75),
	.Q(n_741));
   NAND2_A_OAI21_X2_50_SVT g44481 (.A0N(DPATH_RF_MEMORY_4__9_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN3_n_64),
	.Q(n_740));
   NAND2_A_OAI21_X2_50_SVT g44482 (.A0N(DPATH_RF_MEMORY_18__29_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN76_n_75),
	.Q(n_739));
   NAND2_A_OAI21_X2_50_SVT g44483 (.A0N(DPATH_RF_MEMORY_4__10_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN105_n_134),
	.B1(FE_OFN3_n_64),
	.Q(n_738));
   NAND2_A_OAI21_X2_50_SVT g44484 (.A0N(DPATH_RF_MEMORY_18__30_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN76_n_75),
	.Q(n_737));
   NAND2_A_OAI21_X2_50_SVT g44485 (.A0N(DPATH_RF_MEMORY_18__31_),
	.A1N(FE_OFN76_n_75),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN76_n_75),
	.Q(n_736));
   NAND2_A_OAI21_X2_50_SVT g44486 (.A0N(DPATH_RF_MEMORY_4__11_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN3_n_64),
	.Q(n_735));
   NAND2_A_OAI21_X2_50_SVT g44487 (.A0N(DPATH_RF_MEMORY_4__12_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN3_n_64),
	.Q(n_734));
   NAND2_A_OAI21_X2_50_SVT g44488 (.A0N(DPATH_RF_MEMORY_4__13_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN110_n_142),
	.B1(FE_OFN3_n_64),
	.Q(n_733));
   NAND2_A_OAI21_X2_50_SVT g44489 (.A0N(DPATH_RF_MEMORY_4__14_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN3_n_64),
	.Q(n_732));
   NAND2_A_OAI21_X2_50_SVT g44490 (.A0N(DPATH_RF_MEMORY_4__15_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN3_n_64),
	.Q(n_731));
   NAND2_A_OAI21_X2_50_SVT g44491 (.A0N(DPATH_RF_MEMORY_4__16_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN3_n_64),
	.Q(n_730));
   NAND2_A_OAI21_X2_50_SVT g44492 (.A0N(DPATH_RF_MEMORY_4__19_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN3_n_64),
	.Q(n_729));
   NAND2_A_OAI21_X2_50_SVT g44493 (.A0N(DPATH_RF_MEMORY_4__17_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN3_n_64),
	.Q(n_728));
   NAND2_A_OAI21_X2_50_SVT g44494 (.A0N(DPATH_RF_MEMORY_4__18_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN3_n_64),
	.Q(n_727));
   NAND2_A_OAI21_X2_50_SVT g44495 (.A0N(DPATH_RF_MEMORY_4__20_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN3_n_64),
	.Q(n_726));
   NAND2_A_OAI21_X2_50_SVT g44496 (.A0N(DPATH_RF_MEMORY_4__21_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN3_n_64),
	.Q(n_725));
   NAND2_A_OAI21_X2_50_SVT g44497 (.A0N(DPATH_RF_MEMORY_4__22_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN3_n_64),
	.Q(n_724));
   NAND2_A_OAI21_X2_50_SVT g44498 (.A0N(DPATH_RF_MEMORY_28__8_),
	.A1N(FE_OFN80_n_85),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN80_n_85),
	.Q(n_723));
   NAND2_A_OAI21_X2_50_SVT g44499 (.A0N(DPATH_RF_MEMORY_4__23_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN3_n_64),
	.Q(n_722));
   NAND2_A_OAI21_X2_50_SVT g44500 (.A0N(DPATH_RF_MEMORY_4__24_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN3_n_64),
	.Q(n_721));
   NAND2_A_OAI21_X2_50_SVT g44501 (.A0N(DPATH_RF_MEMORY_4__25_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN3_n_64),
	.Q(n_720));
   NAND2_A_OAI21_X2_50_SVT g44502 (.A0N(DPATH_RF_MEMORY_4__26_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN3_n_64),
	.Q(n_719));
   NAND2_A_OAI21_X2_50_SVT g44503 (.A0N(DPATH_RF_MEMORY_4__27_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN3_n_64),
	.Q(n_718));
   NAND2_A_OAI21_X2_50_SVT g44504 (.A0N(DPATH_RF_MEMORY_20__0_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN93_n_117),
	.B1(FE_OFN77_n_76),
	.Q(n_717));
   NAND2_A_OAI21_X2_50_SVT g44505 (.A0N(DPATH_RF_MEMORY_20__1_),
	.A1N(n_76),
	.B0(FE_OFN108_n_140),
	.B1(n_76),
	.Q(n_716));
   NAND2_A_OAI21_X2_50_SVT g44506 (.A0N(DPATH_RF_MEMORY_4__28_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN3_n_64),
	.Q(n_715));
   NAND2_A_OAI21_X2_50_SVT g44507 (.A0N(DPATH_RF_MEMORY_20__3_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN111_n_144),
	.B1(FE_OFN77_n_76),
	.Q(n_714));
   NAND2_A_OAI21_X2_50_SVT g44508 (.A0N(DPATH_RF_MEMORY_20__4_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN82_n_93),
	.B1(FE_OFN77_n_76),
	.Q(n_713));
   NAND2_A_OAI21_X2_50_SVT g44509 (.A0N(DPATH_RF_MEMORY_4__29_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN3_n_64),
	.Q(n_712));
   NAND2_A_OAI21_X2_50_SVT g44510 (.A0N(DPATH_RF_MEMORY_20__5_),
	.A1N(n_76),
	.B0(FE_OFN116_n_152),
	.B1(n_76),
	.Q(n_711));
   NAND2_A_OAI21_X2_50_SVT g44511 (.A0N(DPATH_RF_MEMORY_4__30_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN3_n_64),
	.Q(n_710));
   NAND2_A_OAI21_X2_50_SVT g44512 (.A0N(DPATH_RF_MEMORY_20__6_),
	.A1N(n_76),
	.B0(FE_OFN107_n_138),
	.B1(n_76),
	.Q(n_709));
   NAND2_A_OAI21_X2_50_SVT g44513 (.A0N(DPATH_RF_MEMORY_4__31_),
	.A1N(FE_OFN3_n_64),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN3_n_64),
	.Q(n_708));
   NAND2_A_OAI21_X2_50_SVT g44514 (.A0N(DPATH_RF_MEMORY_20__7_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN88_n_107),
	.B1(FE_OFN77_n_76),
	.Q(n_707));
   NAND2_A_OAI21_X2_50_SVT g44515 (.A0N(DPATH_RF_MEMORY_20__8_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN106_n_136),
	.B1(FE_OFN77_n_76),
	.Q(n_706));
   NAND2_A_OAI21_X2_50_SVT g44516 (.A0N(DPATH_RF_MEMORY_20__9_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN96_n_121),
	.B1(FE_OFN77_n_76),
	.Q(n_705));
   NAND2_A_OAI21_X2_50_SVT g44517 (.A0N(DPATH_RF_MEMORY_20__10_),
	.A1N(n_76),
	.B0(FE_OFN105_n_134),
	.B1(n_76),
	.Q(n_704));
   NAND2_A_OAI21_X2_50_SVT g44518 (.A0N(DPATH_RF_MEMORY_28__4_),
	.A1N(n_85),
	.B0(FE_OFN82_n_93),
	.B1(n_85),
	.Q(n_703));
   NAND2_A_OAI21_X2_50_SVT g44519 (.A0N(DPATH_RF_MEMORY_20__11_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN103_n_132),
	.B1(FE_OFN77_n_76),
	.Q(n_702));
   NAND2_A_OAI21_X2_50_SVT g44520 (.A0N(DPATH_RF_MEMORY_20__12_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN102_n_130),
	.B1(FE_OFN77_n_76),
	.Q(n_701));
   NAND2_A_OAI21_X2_50_SVT g44521 (.A0N(DPATH_RF_MEMORY_20__13_),
	.A1N(n_76),
	.B0(FE_OFN110_n_142),
	.B1(n_76),
	.Q(n_700));
   NAND2_A_OAI21_X2_50_SVT g44522 (.A0N(DPATH_RF_MEMORY_20__14_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN100_n_127),
	.B1(FE_OFN77_n_76),
	.Q(n_699));
   NAND2_A_OAI21_X2_50_SVT g44523 (.A0N(DPATH_RF_MEMORY_20__15_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN99_n_125),
	.B1(FE_OFN77_n_76),
	.Q(n_698));
   NAND2_A_OAI21_X2_50_SVT g44524 (.A0N(DPATH_RF_MEMORY_20__16_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN117_n_154),
	.B1(FE_OFN77_n_76),
	.Q(n_697));
   NAND2_A_OAI21_X2_50_SVT g44525 (.A0N(DPATH_RF_MEMORY_20__17_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN95_n_119),
	.B1(FE_OFN77_n_76),
	.Q(n_696));
   NAND2_A_OAI21_X2_50_SVT g44526 (.A0N(DPATH_RF_MEMORY_20__18_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN113_n_148),
	.B1(FE_OFN77_n_76),
	.Q(n_695));
   NAND2_A_OAI21_X2_50_SVT g44527 (.A0N(DPATH_RF_MEMORY_20__19_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN92_n_115),
	.B1(FE_OFN77_n_76),
	.Q(n_694));
   NAND2_A_OAI21_X2_50_SVT g44528 (.A0N(DPATH_RF_MEMORY_20__20_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN91_n_113),
	.B1(FE_OFN77_n_76),
	.Q(n_693));
   NAND2_A_OAI21_X2_50_SVT g44529 (.A0N(DPATH_RF_MEMORY_20__21_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN112_n_146),
	.B1(FE_OFN77_n_76),
	.Q(n_692));
   NAND2_A_OAI21_X2_50_SVT g44530 (.A0N(DPATH_RF_MEMORY_20__22_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN114_n_150),
	.B1(FE_OFN77_n_76),
	.Q(n_691));
   NAND2_A_OAI21_X2_50_SVT g44531 (.A0N(DPATH_RF_MEMORY_20__23_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN97_n_123),
	.B1(FE_OFN77_n_76),
	.Q(n_690));
   NAND2_A_OAI21_X2_50_SVT g44532 (.A0N(DPATH_RF_MEMORY_20__24_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN90_n_111),
	.B1(FE_OFN77_n_76),
	.Q(n_689));
   NAND2_A_OAI21_X2_50_SVT g44533 (.A0N(DPATH_RF_MEMORY_20__25_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN89_n_109),
	.B1(FE_OFN77_n_76),
	.Q(n_688));
   NAND2_A_OAI21_X2_50_SVT g44534 (.A0N(DPATH_RF_MEMORY_20__26_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN87_n_105),
	.B1(FE_OFN77_n_76),
	.Q(n_687));
   NAND2_A_OAI21_X2_50_SVT g44535 (.A0N(DPATH_RF_MEMORY_20__27_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN86_n_103),
	.B1(FE_OFN77_n_76),
	.Q(n_686));
   NAND2_A_OAI21_X2_50_SVT g44536 (.A0N(DPATH_RF_MEMORY_20__28_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN85_n_101),
	.B1(FE_OFN77_n_76),
	.Q(n_685));
   NAND2_A_OAI21_X2_50_SVT g44537 (.A0N(DPATH_RF_MEMORY_20__29_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN84_n_99),
	.B1(FE_OFN77_n_76),
	.Q(n_684));
   NAND2_A_OAI21_X2_50_SVT g44538 (.A0N(DPATH_RF_MEMORY_20__30_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN83_n_97),
	.B1(FE_OFN77_n_76),
	.Q(n_683));
   NAND2_A_OAI21_X2_50_SVT g44539 (.A0N(DPATH_RF_MEMORY_20__31_),
	.A1N(FE_OFN77_n_76),
	.B0(FE_OFN119_n_95),
	.B1(FE_OFN77_n_76),
	.Q(n_682));
   MUX2_X2_50_SVT g44540 (.A(DPATH_RF_MEMORY_6__0_),
	.B(n_116),
	.Q(n_681),
	.S0(n_65));
   MUX2_X2_50_SVT g44541 (.A(DPATH_RF_MEMORY_6__1_),
	.B(n_139),
	.Q(n_680),
	.S0(n_65));
   MUX2_X2_50_SVT g44542 (.A(DPATH_RF_MEMORY_6__3_),
	.B(n_143),
	.Q(n_679),
	.S0(n_65));
   MUX2_X2_50_SVT g44543 (.A(DPATH_RF_MEMORY_6__4_),
	.B(n_92),
	.Q(n_678),
	.S0(n_65));
   MUX2_X2_50_SVT g44544 (.A(DPATH_RF_MEMORY_6__5_),
	.B(n_151),
	.Q(n_677),
	.S0(n_65));
   MUX2_X2_50_SVT g44545 (.A(DPATH_RF_MEMORY_6__6_),
	.B(n_137),
	.Q(n_676),
	.S0(n_65));
   MUX2_X2_50_SVT g44546 (.A(DPATH_RF_MEMORY_6__7_),
	.B(n_106),
	.Q(n_675),
	.S0(n_65));
   MUX2_X2_50_SVT g44547 (.A(DPATH_RF_MEMORY_6__8_),
	.B(n_135),
	.Q(n_674),
	.S0(n_65));
   MUX2_X2_50_SVT g44548 (.A(DPATH_RF_MEMORY_6__9_),
	.B(n_120),
	.Q(n_673),
	.S0(n_65));
   MUX2_X2_50_SVT g44549 (.A(DPATH_RF_MEMORY_6__10_),
	.B(n_133),
	.Q(n_672),
	.S0(n_65));
   MUX2_X2_50_SVT g44550 (.A(DPATH_RF_MEMORY_6__11_),
	.B(n_131),
	.Q(n_671),
	.S0(n_65));
   MUX2_X2_50_SVT g44551 (.A(DPATH_RF_MEMORY_6__12_),
	.B(n_129),
	.Q(n_670),
	.S0(n_65));
   MUX2_X2_50_SVT g44552 (.A(DPATH_RF_MEMORY_6__13_),
	.B(n_141),
	.Q(n_669),
	.S0(n_65));
   MUX2_X2_50_SVT g44553 (.A(DPATH_RF_MEMORY_6__14_),
	.B(n_126),
	.Q(n_668),
	.S0(n_65));
   MUX2_X2_50_SVT g44554 (.A(DPATH_RF_MEMORY_6__15_),
	.B(n_124),
	.Q(n_667),
	.S0(n_65));
   MUX2_X2_50_SVT g44555 (.A(DPATH_RF_MEMORY_6__18_),
	.B(n_147),
	.Q(n_666),
	.S0(n_65));
   MUX2_X2_50_SVT g44556 (.A(DPATH_RF_MEMORY_6__16_),
	.B(n_153),
	.Q(n_665),
	.S0(n_65));
   MUX2_X2_50_SVT g44557 (.A(DPATH_RF_MEMORY_6__17_),
	.B(n_118),
	.Q(n_664),
	.S0(n_65));
   MUX2_X2_50_SVT g44558 (.A(DPATH_RF_MEMORY_6__19_),
	.B(n_114),
	.Q(n_663),
	.S0(n_65));
   MUX2_X2_50_SVT g44559 (.A(DPATH_RF_MEMORY_6__20_),
	.B(n_112),
	.Q(n_662),
	.S0(n_65));
   MUX2_X2_50_SVT g44560 (.A(DPATH_RF_MEMORY_6__21_),
	.B(n_145),
	.Q(n_661),
	.S0(n_65));
   MUX2_X2_50_SVT g44561 (.A(DPATH_RF_MEMORY_6__22_),
	.B(n_149),
	.Q(n_660),
	.S0(n_65));
   MUX2_X2_50_SVT g44562 (.A(DPATH_RF_MEMORY_6__23_),
	.B(n_122),
	.Q(n_659),
	.S0(n_65));
   MUX2_X2_50_SVT g44563 (.A(DPATH_RF_MEMORY_6__24_),
	.B(n_110),
	.Q(n_658),
	.S0(n_65));
   MUX2_X2_50_SVT g44564 (.A(DPATH_RF_MEMORY_6__25_),
	.B(n_108),
	.Q(n_657),
	.S0(n_65));
   MUX2_X2_50_SVT g44565 (.A(DPATH_RF_MEMORY_6__26_),
	.B(n_104),
	.Q(n_656),
	.S0(n_65));
   MUX2_X2_50_SVT g44566 (.A(DPATH_RF_MEMORY_6__27_),
	.B(n_102),
	.Q(n_655),
	.S0(n_65));
   MUX2_X2_50_SVT g44567 (.A(DPATH_RF_MEMORY_6__28_),
	.B(n_100),
	.Q(n_654),
	.S0(n_65));
   MUX2_X2_50_SVT g44568 (.A(DPATH_RF_MEMORY_6__29_),
	.B(n_98),
	.Q(n_653),
	.S0(n_65));
   MUX2_X2_50_SVT g44569 (.A(DPATH_RF_MEMORY_6__30_),
	.B(n_96),
	.Q(n_652),
	.S0(n_65));
   MUX2_X2_50_SVT g44570 (.A(DPATH_RF_MEMORY_6__31_),
	.B(n_94),
	.Q(n_651),
	.S0(n_65));
   MUX2_X2_50_SVT g44571 (.A(DPATH_RF_MEMORY_27__0_),
	.B(n_116),
	.Q(n_650),
	.S0(n_66));
   MUX2_X2_50_SVT g44572 (.A(DPATH_RF_MEMORY_27__1_),
	.B(n_139),
	.Q(n_649),
	.S0(n_66));
   MUX2_X2_50_SVT g44573 (.A(DPATH_RF_MEMORY_27__3_),
	.B(n_143),
	.Q(n_648),
	.S0(n_66));
   MUX2_X2_50_SVT g44574 (.A(DPATH_RF_MEMORY_27__4_),
	.B(n_92),
	.Q(n_647),
	.S0(n_66));
   MUX2_X2_50_SVT g44575 (.A(DPATH_RF_MEMORY_27__5_),
	.B(n_151),
	.Q(n_646),
	.S0(n_66));
   MUX2_X2_50_SVT g44576 (.A(DPATH_RF_MEMORY_27__6_),
	.B(n_137),
	.Q(n_645),
	.S0(n_66));
   MUX2_X2_50_SVT g44577 (.A(DPATH_RF_MEMORY_27__7_),
	.B(n_106),
	.Q(n_644),
	.S0(n_66));
   MUX2_X2_50_SVT g44578 (.A(DPATH_RF_MEMORY_27__8_),
	.B(n_135),
	.Q(n_643),
	.S0(n_66));
   MUX2_X2_50_SVT g44579 (.A(DPATH_RF_MEMORY_27__9_),
	.B(n_120),
	.Q(n_642),
	.S0(n_66));
   MUX2_X2_50_SVT g44580 (.A(DPATH_RF_MEMORY_27__10_),
	.B(n_133),
	.Q(n_641),
	.S0(n_66));
   MUX2_X2_50_SVT g44581 (.A(DPATH_RF_MEMORY_27__11_),
	.B(n_131),
	.Q(n_640),
	.S0(n_66));
   MUX2_X2_50_SVT g44582 (.A(DPATH_RF_MEMORY_27__12_),
	.B(n_129),
	.Q(n_639),
	.S0(n_66));
   MUX2_X2_50_SVT g44583 (.A(DPATH_RF_MEMORY_27__13_),
	.B(n_141),
	.Q(n_638),
	.S0(n_66));
   MUX2_X2_50_SVT g44584 (.A(DPATH_RF_MEMORY_27__14_),
	.B(n_126),
	.Q(n_637),
	.S0(n_66));
   MUX2_X2_50_SVT g44585 (.A(DPATH_RF_MEMORY_27__15_),
	.B(n_124),
	.Q(n_636),
	.S0(n_66));
   MUX2_X2_50_SVT g44586 (.A(DPATH_RF_MEMORY_27__16_),
	.B(n_153),
	.Q(n_635),
	.S0(n_66));
   MUX2_X2_50_SVT g44587 (.A(DPATH_RF_MEMORY_27__17_),
	.B(n_118),
	.Q(n_634),
	.S0(n_66));
   MUX2_X2_50_SVT g44588 (.A(DPATH_RF_MEMORY_27__18_),
	.B(n_147),
	.Q(n_633),
	.S0(n_66));
   MUX2_X2_50_SVT g44589 (.A(DPATH_RF_MEMORY_27__19_),
	.B(n_114),
	.Q(n_632),
	.S0(n_66));
   MUX2_X2_50_SVT g44590 (.A(DPATH_RF_MEMORY_27__20_),
	.B(n_112),
	.Q(n_631),
	.S0(n_66));
   MUX2_X2_50_SVT g44591 (.A(DPATH_RF_MEMORY_27__21_),
	.B(n_145),
	.Q(n_630),
	.S0(n_66));
   MUX2_X2_50_SVT g44592 (.A(DPATH_RF_MEMORY_27__22_),
	.B(n_149),
	.Q(n_629),
	.S0(n_66));
   MUX2_X2_50_SVT g44593 (.A(DPATH_RF_MEMORY_27__23_),
	.B(n_122),
	.Q(n_628),
	.S0(n_66));
   MUX2_X2_50_SVT g44594 (.A(DPATH_RF_MEMORY_27__24_),
	.B(n_110),
	.Q(n_627),
	.S0(n_66));
   MUX2_X2_50_SVT g44595 (.A(DPATH_RF_MEMORY_27__25_),
	.B(n_108),
	.Q(n_626),
	.S0(n_66));
   MUX2_X2_50_SVT g44596 (.A(DPATH_RF_MEMORY_27__26_),
	.B(n_104),
	.Q(n_625),
	.S0(n_66));
   MUX2_X2_50_SVT g44597 (.A(DPATH_RF_MEMORY_27__27_),
	.B(n_102),
	.Q(n_624),
	.S0(n_66));
   MUX2_X2_50_SVT g44598 (.A(DPATH_RF_MEMORY_27__28_),
	.B(n_100),
	.Q(n_623),
	.S0(n_66));
   MUX2_X2_50_SVT g44599 (.A(DPATH_RF_MEMORY_27__29_),
	.B(n_98),
	.Q(n_622),
	.S0(n_66));
   MUX2_X2_50_SVT g44600 (.A(DPATH_RF_MEMORY_27__30_),
	.B(n_96),
	.Q(n_621),
	.S0(n_66));
   MUX2_X2_50_SVT g44601 (.A(DPATH_RF_MEMORY_27__31_),
	.B(n_94),
	.Q(n_620),
	.S0(n_66));
   MUX2_X2_50_SVT g44602 (.A(DPATH_RF_MEMORY_31__0_),
	.B(n_116),
	.Q(n_619),
	.S0(n_68));
   MUX2_X2_50_SVT g44603 (.A(DPATH_RF_MEMORY_31__1_),
	.B(n_139),
	.Q(n_618),
	.S0(n_68));
   MUX2_X2_50_SVT g44604 (.A(DPATH_RF_MEMORY_31__3_),
	.B(n_143),
	.Q(n_617),
	.S0(n_68));
   MUX2_X2_50_SVT g44605 (.A(DPATH_RF_MEMORY_31__4_),
	.B(n_92),
	.Q(n_616),
	.S0(n_68));
   MUX2_X2_50_SVT g44606 (.A(DPATH_RF_MEMORY_31__5_),
	.B(n_151),
	.Q(n_615),
	.S0(n_68));
   MUX2_X2_50_SVT g44607 (.A(DPATH_RF_MEMORY_31__6_),
	.B(n_137),
	.Q(n_614),
	.S0(n_68));
   MUX2_X2_50_SVT g44608 (.A(DPATH_RF_MEMORY_31__7_),
	.B(n_106),
	.Q(n_613),
	.S0(n_68));
   MUX2_X2_50_SVT g44609 (.A(DPATH_RF_MEMORY_31__8_),
	.B(n_135),
	.Q(n_612),
	.S0(n_68));
   MUX2_X2_50_SVT g44610 (.A(DPATH_RF_MEMORY_31__9_),
	.B(n_120),
	.Q(n_611),
	.S0(n_68));
   MUX2_X2_50_SVT g44611 (.A(DPATH_RF_MEMORY_31__10_),
	.B(n_133),
	.Q(n_610),
	.S0(n_68));
   MUX2_X2_50_SVT g44612 (.A(DPATH_RF_MEMORY_31__11_),
	.B(n_131),
	.Q(n_609),
	.S0(n_68));
   MUX2_X2_50_SVT g44613 (.A(DPATH_RF_MEMORY_31__12_),
	.B(n_129),
	.Q(n_608),
	.S0(n_68));
   MUX2_X2_50_SVT g44614 (.A(DPATH_RF_MEMORY_31__13_),
	.B(n_141),
	.Q(n_607),
	.S0(n_68));
   MUX2_X2_50_SVT g44615 (.A(DPATH_RF_MEMORY_31__14_),
	.B(n_126),
	.Q(n_606),
	.S0(n_68));
   MUX2_X2_50_SVT g44616 (.A(DPATH_RF_MEMORY_31__15_),
	.B(n_124),
	.Q(n_605),
	.S0(n_68));
   MUX2_X2_50_SVT g44617 (.A(DPATH_RF_MEMORY_31__16_),
	.B(n_153),
	.Q(n_604),
	.S0(n_68));
   MUX2_X2_50_SVT g44618 (.A(DPATH_RF_MEMORY_31__17_),
	.B(n_118),
	.Q(n_603),
	.S0(n_68));
   MUX2_X2_50_SVT g44619 (.A(DPATH_RF_MEMORY_31__18_),
	.B(n_147),
	.Q(n_602),
	.S0(n_68));
   MUX2_X2_50_SVT g44620 (.A(DPATH_RF_MEMORY_31__19_),
	.B(n_114),
	.Q(n_601),
	.S0(n_68));
   MUX2_X2_50_SVT g44621 (.A(DPATH_RF_MEMORY_31__20_),
	.B(n_112),
	.Q(n_600),
	.S0(n_68));
   MUX2_X2_50_SVT g44622 (.A(DPATH_RF_MEMORY_31__21_),
	.B(n_145),
	.Q(n_599),
	.S0(n_68));
   MUX2_X2_50_SVT g44623 (.A(DPATH_RF_MEMORY_31__22_),
	.B(n_149),
	.Q(n_598),
	.S0(n_68));
   MUX2_X2_50_SVT g44624 (.A(DPATH_RF_MEMORY_31__23_),
	.B(n_122),
	.Q(n_597),
	.S0(n_68));
   MUX2_X2_50_SVT g44625 (.A(DPATH_RF_MEMORY_31__24_),
	.B(n_110),
	.Q(n_596),
	.S0(n_68));
   MUX2_X2_50_SVT g44626 (.A(DPATH_RF_MEMORY_31__25_),
	.B(n_108),
	.Q(n_595),
	.S0(n_68));
   MUX2_X2_50_SVT g44627 (.A(DPATH_RF_MEMORY_31__26_),
	.B(n_104),
	.Q(n_594),
	.S0(n_68));
   MUX2_X2_50_SVT g44628 (.A(DPATH_RF_MEMORY_31__27_),
	.B(n_102),
	.Q(n_593),
	.S0(n_68));
   MUX2_X2_50_SVT g44629 (.A(DPATH_RF_MEMORY_31__28_),
	.B(n_100),
	.Q(n_592),
	.S0(n_68));
   MUX2_X2_50_SVT g44630 (.A(DPATH_RF_MEMORY_31__29_),
	.B(n_98),
	.Q(n_591),
	.S0(n_68));
   MUX2_X2_50_SVT g44631 (.A(DPATH_RF_MEMORY_31__30_),
	.B(n_96),
	.Q(n_590),
	.S0(n_68));
   MUX2_X2_50_SVT g44632 (.A(DPATH_RF_MEMORY_31__31_),
	.B(n_94),
	.Q(n_589),
	.S0(n_68));
   MUX2_X2_50_SVT g44633 (.A(DPATH_RF_MEMORY_2__0_),
	.B(n_116),
	.Q(n_588),
	.S0(n_63));
   MUX2_X2_50_SVT g44634 (.A(DPATH_RF_MEMORY_2__1_),
	.B(n_139),
	.Q(n_587),
	.S0(n_63));
   MUX2_X2_50_SVT g44635 (.A(DPATH_RF_MEMORY_2__4_),
	.B(n_92),
	.Q(n_586),
	.S0(n_63));
   MUX2_X2_50_SVT g44636 (.A(DPATH_RF_MEMORY_2__3_),
	.B(n_143),
	.Q(n_585),
	.S0(n_63));
   MUX2_X2_50_SVT g44637 (.A(DPATH_RF_MEMORY_2__5_),
	.B(n_151),
	.Q(n_584),
	.S0(n_63));
   MUX2_X2_50_SVT g44638 (.A(DPATH_RF_MEMORY_2__6_),
	.B(n_137),
	.Q(n_583),
	.S0(n_63));
   MUX2_X2_50_SVT g44639 (.A(DPATH_RF_MEMORY_2__7_),
	.B(n_106),
	.Q(n_582),
	.S0(n_63));
   MUX2_X2_50_SVT g44640 (.A(DPATH_RF_MEMORY_2__8_),
	.B(n_135),
	.Q(n_581),
	.S0(n_63));
   MUX2_X2_50_SVT g44641 (.A(DPATH_RF_MEMORY_2__9_),
	.B(n_120),
	.Q(n_580),
	.S0(n_63));
   MUX2_X2_50_SVT g44642 (.A(DPATH_RF_MEMORY_2__10_),
	.B(n_133),
	.Q(n_579),
	.S0(n_63));
   MUX2_X2_50_SVT g44643 (.A(DPATH_RF_MEMORY_2__11_),
	.B(n_131),
	.Q(n_578),
	.S0(n_63));
   MUX2_X2_50_SVT g44644 (.A(DPATH_RF_MEMORY_2__12_),
	.B(n_129),
	.Q(n_577),
	.S0(n_63));
   MUX2_X2_50_SVT g44645 (.A(DPATH_RF_MEMORY_2__13_),
	.B(n_141),
	.Q(n_576),
	.S0(n_63));
   MUX2_X2_50_SVT g44646 (.A(DPATH_RF_MEMORY_2__14_),
	.B(n_126),
	.Q(n_575),
	.S0(n_63));
   MUX2_X2_50_SVT g44647 (.A(DPATH_RF_MEMORY_2__15_),
	.B(n_124),
	.Q(n_574),
	.S0(n_63));
   MUX2_X2_50_SVT g44648 (.A(DPATH_RF_MEMORY_2__16_),
	.B(n_153),
	.Q(n_573),
	.S0(n_63));
   MUX2_X2_50_SVT g44649 (.A(DPATH_RF_MEMORY_2__17_),
	.B(n_118),
	.Q(n_572),
	.S0(n_63));
   MUX2_X2_50_SVT g44650 (.A(DPATH_RF_MEMORY_2__20_),
	.B(n_112),
	.Q(n_571),
	.S0(n_63));
   MUX2_X2_50_SVT g44651 (.A(DPATH_RF_MEMORY_2__18_),
	.B(n_147),
	.Q(n_570),
	.S0(n_63));
   MUX2_X2_50_SVT g44652 (.A(DPATH_RF_MEMORY_2__19_),
	.B(n_114),
	.Q(n_569),
	.S0(n_63));
   MUX2_X2_50_SVT g44653 (.A(DPATH_RF_MEMORY_2__21_),
	.B(n_145),
	.Q(n_568),
	.S0(n_63));
   MUX2_X2_50_SVT g44654 (.A(DPATH_RF_MEMORY_2__22_),
	.B(n_149),
	.Q(n_567),
	.S0(n_63));
   MUX2_X2_50_SVT g44655 (.A(DPATH_RF_MEMORY_2__23_),
	.B(n_122),
	.Q(n_566),
	.S0(n_63));
   MUX2_X2_50_SVT g44656 (.A(DPATH_RF_MEMORY_2__24_),
	.B(n_110),
	.Q(n_565),
	.S0(n_63));
   MUX2_X2_50_SVT g44657 (.A(DPATH_RF_MEMORY_2__25_),
	.B(n_108),
	.Q(n_564),
	.S0(n_63));
   MUX2_X2_50_SVT g44658 (.A(DPATH_RF_MEMORY_2__26_),
	.B(n_104),
	.Q(n_563),
	.S0(n_63));
   MUX2_X2_50_SVT g44659 (.A(DPATH_RF_MEMORY_2__27_),
	.B(n_102),
	.Q(n_562),
	.S0(n_63));
   MUX2_X2_50_SVT g44660 (.A(DPATH_RF_MEMORY_2__28_),
	.B(n_100),
	.Q(n_561),
	.S0(n_63));
   MUX2_X2_50_SVT g44661 (.A(DPATH_RF_MEMORY_2__29_),
	.B(n_98),
	.Q(n_560),
	.S0(n_63));
   MUX2_X2_50_SVT g44662 (.A(DPATH_RF_MEMORY_2__30_),
	.B(n_96),
	.Q(n_559),
	.S0(n_63));
   MUX2_X2_50_SVT g44663 (.A(DPATH_RF_MEMORY_2__31_),
	.B(n_94),
	.Q(n_558),
	.S0(n_63));
   MUX2_X2_50_SVT g44664 (.A(DPATH_RF_MEMORY_5__18_),
	.B(n_147),
	.Q(n_557),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44665 (.A(DPATH_RF_MEMORY_21__11_),
	.B(n_131),
	.Q(n_556),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44666 (.A(DPATH_RF_MEMORY_21__12_),
	.B(n_129),
	.Q(n_555),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44667 (.A(DPATH_RF_MEMORY_21__13_),
	.B(n_141),
	.Q(n_554),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44668 (.A(DPATH_RF_MEMORY_21__14_),
	.B(n_126),
	.Q(n_553),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44669 (.A(DPATH_RF_MEMORY_21__15_),
	.B(n_124),
	.Q(n_552),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44670 (.A(DPATH_RF_MEMORY_5__19_),
	.B(n_114),
	.Q(n_551),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44671 (.A(DPATH_RF_MEMORY_21__16_),
	.B(n_153),
	.Q(n_550),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44672 (.A(DPATH_RF_MEMORY_5__20_),
	.B(n_112),
	.Q(n_549),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44673 (.A(DPATH_RF_MEMORY_21__17_),
	.B(n_118),
	.Q(n_548),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44674 (.A(DPATH_RF_MEMORY_21__18_),
	.B(n_147),
	.Q(n_547),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44675 (.A(DPATH_RF_MEMORY_21__19_),
	.B(n_114),
	.Q(n_546),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44676 (.A(DPATH_RF_MEMORY_5__17_),
	.B(n_118),
	.Q(n_545),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44677 (.A(DPATH_RF_MEMORY_21__20_),
	.B(n_112),
	.Q(n_544),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44678 (.A(DPATH_RF_MEMORY_5__21_),
	.B(n_145),
	.Q(n_543),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44679 (.A(DPATH_RF_MEMORY_21__21_),
	.B(n_145),
	.Q(n_542),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44680 (.A(DPATH_RF_MEMORY_5__22_),
	.B(n_149),
	.Q(n_541),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44681 (.A(DPATH_RF_MEMORY_21__22_),
	.B(n_149),
	.Q(n_540),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44682 (.A(DPATH_RF_MEMORY_5__23_),
	.B(n_122),
	.Q(n_539),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44683 (.A(DPATH_RF_MEMORY_21__23_),
	.B(n_122),
	.Q(n_538),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44684 (.A(DPATH_RF_MEMORY_21__24_),
	.B(n_110),
	.Q(n_537),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44685 (.A(DPATH_RF_MEMORY_21__25_),
	.B(n_108),
	.Q(n_536),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44686 (.A(DPATH_RF_MEMORY_5__24_),
	.B(n_110),
	.Q(n_535),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44687 (.A(DPATH_RF_MEMORY_21__26_),
	.B(n_104),
	.Q(n_534),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44688 (.A(DPATH_RF_MEMORY_21__27_),
	.B(n_102),
	.Q(n_533),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44689 (.A(DPATH_RF_MEMORY_5__25_),
	.B(n_108),
	.Q(n_532),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44690 (.A(DPATH_RF_MEMORY_21__28_),
	.B(n_100),
	.Q(n_531),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44691 (.A(DPATH_RF_MEMORY_5__26_),
	.B(n_104),
	.Q(n_530),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44692 (.A(DPATH_RF_MEMORY_21__29_),
	.B(n_98),
	.Q(n_529),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44693 (.A(DPATH_RF_MEMORY_21__30_),
	.B(n_96),
	.Q(n_528),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44694 (.A(DPATH_RF_MEMORY_5__27_),
	.B(n_102),
	.Q(n_527),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44695 (.A(DPATH_RF_MEMORY_21__31_),
	.B(n_94),
	.Q(n_526),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44696 (.A(DPATH_RF_MEMORY_5__28_),
	.B(n_100),
	.Q(n_525),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44697 (.A(DPATH_RF_MEMORY_5__29_),
	.B(n_98),
	.Q(n_524),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44698 (.A(DPATH_RF_MEMORY_5__30_),
	.B(n_96),
	.Q(n_523),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44699 (.A(DPATH_RF_MEMORY_5__31_),
	.B(n_94),
	.Q(n_522),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44700 (.A(DPATH_RF_MEMORY_13__0_),
	.B(n_116),
	.Q(n_521),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44701 (.A(DPATH_RF_MEMORY_13__1_),
	.B(n_139),
	.Q(n_520),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44702 (.A(DPATH_RF_MEMORY_13__3_),
	.B(n_143),
	.Q(n_519),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44703 (.A(DPATH_RF_MEMORY_13__4_),
	.B(n_92),
	.Q(n_518),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44704 (.A(DPATH_RF_MEMORY_13__5_),
	.B(n_151),
	.Q(n_517),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44705 (.A(DPATH_RF_MEMORY_13__6_),
	.B(n_137),
	.Q(n_516),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44706 (.A(DPATH_RF_MEMORY_13__7_),
	.B(n_106),
	.Q(n_515),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44707 (.A(DPATH_RF_MEMORY_13__8_),
	.B(n_135),
	.Q(n_514),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44708 (.A(DPATH_RF_MEMORY_13__9_),
	.B(n_120),
	.Q(n_513),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44709 (.A(DPATH_RF_MEMORY_13__10_),
	.B(n_133),
	.Q(n_512),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44710 (.A(DPATH_RF_MEMORY_13__11_),
	.B(n_131),
	.Q(n_511),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44711 (.A(DPATH_RF_MEMORY_13__12_),
	.B(n_129),
	.Q(n_510),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44712 (.A(DPATH_RF_MEMORY_13__13_),
	.B(n_141),
	.Q(n_509),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44713 (.A(DPATH_RF_MEMORY_13__15_),
	.B(n_124),
	.Q(n_508),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44714 (.A(DPATH_RF_MEMORY_13__16_),
	.B(n_153),
	.Q(n_507),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44715 (.A(DPATH_RF_MEMORY_13__14_),
	.B(n_126),
	.Q(n_506),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44716 (.A(DPATH_RF_MEMORY_13__17_),
	.B(n_118),
	.Q(n_505),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44717 (.A(DPATH_RF_MEMORY_13__18_),
	.B(n_147),
	.Q(n_504),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44718 (.A(DPATH_RF_MEMORY_13__19_),
	.B(n_114),
	.Q(n_503),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44719 (.A(DPATH_RF_MEMORY_13__20_),
	.B(n_112),
	.Q(n_502),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44720 (.A(DPATH_RF_MEMORY_13__21_),
	.B(n_145),
	.Q(n_501),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44721 (.A(DPATH_RF_MEMORY_13__22_),
	.B(n_149),
	.Q(n_500),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44722 (.A(DPATH_RF_MEMORY_13__23_),
	.B(n_122),
	.Q(n_499),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44723 (.A(DPATH_RF_MEMORY_13__24_),
	.B(n_110),
	.Q(n_498),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44724 (.A(DPATH_RF_MEMORY_13__25_),
	.B(n_108),
	.Q(n_497),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44725 (.A(DPATH_RF_MEMORY_13__26_),
	.B(n_104),
	.Q(n_496),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44726 (.A(DPATH_RF_MEMORY_13__27_),
	.B(n_102),
	.Q(n_495),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44727 (.A(DPATH_RF_MEMORY_13__28_),
	.B(n_100),
	.Q(n_494),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44728 (.A(DPATH_RF_MEMORY_13__29_),
	.B(n_98),
	.Q(n_493),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44729 (.A(DPATH_RF_MEMORY_13__30_),
	.B(n_96),
	.Q(n_492),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44730 (.A(DPATH_RF_MEMORY_13__31_),
	.B(n_94),
	.Q(n_491),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g44731 (.A(DPATH_RF_MEMORY_5__0_),
	.B(n_116),
	.Q(n_490),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44732 (.A(DPATH_RF_MEMORY_5__3_),
	.B(n_143),
	.Q(n_489),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44733 (.A(DPATH_RF_MEMORY_5__1_),
	.B(n_139),
	.Q(n_488),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44734 (.A(DPATH_RF_MEMORY_5__4_),
	.B(n_92),
	.Q(n_487),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44735 (.A(DPATH_RF_MEMORY_5__5_),
	.B(n_151),
	.Q(n_486),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44736 (.A(DPATH_RF_MEMORY_5__6_),
	.B(n_137),
	.Q(n_485),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44737 (.A(DPATH_RF_MEMORY_5__7_),
	.B(n_106),
	.Q(n_484),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44738 (.A(DPATH_RF_MEMORY_5__8_),
	.B(n_135),
	.Q(n_483),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44739 (.A(DPATH_RF_MEMORY_5__9_),
	.B(n_120),
	.Q(n_482),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44740 (.A(DPATH_RF_MEMORY_5__10_),
	.B(n_133),
	.Q(n_481),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44741 (.A(DPATH_RF_MEMORY_5__11_),
	.B(n_131),
	.Q(n_480),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44742 (.A(DPATH_RF_MEMORY_21__0_),
	.B(n_116),
	.Q(n_479),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44743 (.A(DPATH_RF_MEMORY_21__1_),
	.B(n_139),
	.Q(n_478),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44744 (.A(DPATH_RF_MEMORY_5__12_),
	.B(n_129),
	.Q(n_477),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44745 (.A(DPATH_RF_MEMORY_21__3_),
	.B(n_143),
	.Q(n_476),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44746 (.A(DPATH_RF_MEMORY_21__4_),
	.B(n_92),
	.Q(n_475),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44747 (.A(DPATH_RF_MEMORY_5__13_),
	.B(n_141),
	.Q(n_474),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44748 (.A(DPATH_RF_MEMORY_21__5_),
	.B(n_151),
	.Q(n_473),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44749 (.A(DPATH_RF_MEMORY_5__14_),
	.B(n_126),
	.Q(n_472),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44750 (.A(DPATH_RF_MEMORY_21__6_),
	.B(n_137),
	.Q(n_471),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44751 (.A(DPATH_RF_MEMORY_5__15_),
	.B(n_124),
	.Q(n_470),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44752 (.A(DPATH_RF_MEMORY_21__7_),
	.B(n_106),
	.Q(n_469),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44753 (.A(DPATH_RF_MEMORY_21__8_),
	.B(n_135),
	.Q(n_468),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44754 (.A(DPATH_RF_MEMORY_21__9_),
	.B(n_120),
	.Q(n_467),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44755 (.A(DPATH_RF_MEMORY_5__16_),
	.B(n_153),
	.Q(n_466),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g44756 (.A(DPATH_RF_MEMORY_21__10_),
	.B(n_133),
	.Q(n_465),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g44757 (.A(DPATH_RF_MEMORY_23__0_),
	.B(n_116),
	.Q(n_464),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44758 (.A(DPATH_RF_MEMORY_23__1_),
	.B(n_139),
	.Q(n_463),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44759 (.A(DPATH_RF_MEMORY_23__3_),
	.B(n_143),
	.Q(n_462),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44760 (.A(DPATH_RF_MEMORY_23__4_),
	.B(n_92),
	.Q(n_461),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44761 (.A(DPATH_RF_MEMORY_23__5_),
	.B(n_151),
	.Q(n_460),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44762 (.A(DPATH_RF_MEMORY_23__6_),
	.B(n_137),
	.Q(n_459),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44763 (.A(DPATH_RF_MEMORY_23__7_),
	.B(n_106),
	.Q(n_458),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44764 (.A(DPATH_RF_MEMORY_23__8_),
	.B(n_135),
	.Q(n_457),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44765 (.A(DPATH_RF_MEMORY_23__9_),
	.B(n_120),
	.Q(n_456),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44766 (.A(DPATH_RF_MEMORY_23__10_),
	.B(n_133),
	.Q(n_455),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44767 (.A(DPATH_RF_MEMORY_23__11_),
	.B(n_131),
	.Q(n_454),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44768 (.A(DPATH_RF_MEMORY_23__12_),
	.B(n_129),
	.Q(n_453),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44769 (.A(DPATH_RF_MEMORY_23__13_),
	.B(n_141),
	.Q(n_452),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44770 (.A(DPATH_RF_MEMORY_23__14_),
	.B(n_126),
	.Q(n_451),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44771 (.A(DPATH_RF_MEMORY_23__15_),
	.B(n_124),
	.Q(n_450),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44772 (.A(DPATH_RF_MEMORY_23__16_),
	.B(n_153),
	.Q(n_449),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44773 (.A(DPATH_RF_MEMORY_23__17_),
	.B(n_118),
	.Q(n_448),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44774 (.A(DPATH_RF_MEMORY_23__18_),
	.B(n_147),
	.Q(n_447),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44775 (.A(DPATH_RF_MEMORY_23__19_),
	.B(n_114),
	.Q(n_446),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44776 (.A(DPATH_RF_MEMORY_23__20_),
	.B(n_112),
	.Q(n_445),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44777 (.A(DPATH_RF_MEMORY_23__21_),
	.B(n_145),
	.Q(n_444),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44778 (.A(DPATH_RF_MEMORY_23__22_),
	.B(n_149),
	.Q(n_443),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44779 (.A(DPATH_RF_MEMORY_23__23_),
	.B(n_122),
	.Q(n_442),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44780 (.A(DPATH_RF_MEMORY_23__24_),
	.B(n_110),
	.Q(n_441),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44781 (.A(DPATH_RF_MEMORY_23__25_),
	.B(n_108),
	.Q(n_440),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44782 (.A(DPATH_RF_MEMORY_23__26_),
	.B(n_104),
	.Q(n_439),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44783 (.A(DPATH_RF_MEMORY_23__27_),
	.B(n_102),
	.Q(n_438),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44784 (.A(DPATH_RF_MEMORY_23__28_),
	.B(n_100),
	.Q(n_437),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44785 (.A(DPATH_RF_MEMORY_23__29_),
	.B(n_98),
	.Q(n_436),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44786 (.A(DPATH_RF_MEMORY_23__30_),
	.B(n_96),
	.Q(n_435),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44787 (.A(DPATH_RF_MEMORY_23__31_),
	.B(n_94),
	.Q(n_434),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g44788 (.A(DPATH_RF_MEMORY_7__0_),
	.B(n_116),
	.Q(n_433),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44789 (.A(DPATH_RF_MEMORY_7__3_),
	.B(n_143),
	.Q(n_432),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44790 (.A(DPATH_RF_MEMORY_7__1_),
	.B(n_139),
	.Q(n_431),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44791 (.A(DPATH_RF_MEMORY_7__5_),
	.B(n_151),
	.Q(n_430),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44792 (.A(DPATH_RF_MEMORY_7__4_),
	.B(n_92),
	.Q(n_429),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44793 (.A(DPATH_RF_MEMORY_7__6_),
	.B(n_137),
	.Q(n_428),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44794 (.A(DPATH_RF_MEMORY_7__7_),
	.B(n_106),
	.Q(n_427),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44795 (.A(DPATH_RF_MEMORY_7__8_),
	.B(n_135),
	.Q(n_426),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44796 (.A(DPATH_RF_MEMORY_7__9_),
	.B(n_120),
	.Q(n_425),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44797 (.A(DPATH_RF_MEMORY_7__10_),
	.B(n_133),
	.Q(n_424),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44798 (.A(DPATH_RF_MEMORY_7__11_),
	.B(n_131),
	.Q(n_423),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44799 (.A(DPATH_RF_MEMORY_7__13_),
	.B(n_141),
	.Q(n_422),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44800 (.A(DPATH_RF_MEMORY_7__12_),
	.B(n_129),
	.Q(n_421),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44801 (.A(DPATH_RF_MEMORY_7__14_),
	.B(n_126),
	.Q(n_420),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44802 (.A(DPATH_RF_MEMORY_7__15_),
	.B(n_124),
	.Q(n_419),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44803 (.A(DPATH_RF_MEMORY_7__16_),
	.B(n_153),
	.Q(n_418),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44804 (.A(DPATH_RF_MEMORY_7__17_),
	.B(n_118),
	.Q(n_417),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44805 (.A(DPATH_RF_MEMORY_7__19_),
	.B(n_114),
	.Q(n_416),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44806 (.A(DPATH_RF_MEMORY_7__18_),
	.B(n_147),
	.Q(n_415),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44807 (.A(DPATH_RF_MEMORY_7__21_),
	.B(n_145),
	.Q(n_414),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44808 (.A(DPATH_RF_MEMORY_7__20_),
	.B(n_112),
	.Q(n_413),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44809 (.A(DPATH_RF_MEMORY_7__22_),
	.B(n_149),
	.Q(n_412),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44810 (.A(DPATH_RF_MEMORY_7__23_),
	.B(n_122),
	.Q(n_411),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44811 (.A(DPATH_RF_MEMORY_7__24_),
	.B(n_110),
	.Q(n_410),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44812 (.A(DPATH_RF_MEMORY_7__25_),
	.B(n_108),
	.Q(n_409),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44813 (.A(DPATH_RF_MEMORY_7__26_),
	.B(n_104),
	.Q(n_408),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44814 (.A(DPATH_RF_MEMORY_7__27_),
	.B(n_102),
	.Q(n_407),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44815 (.A(DPATH_RF_MEMORY_7__28_),
	.B(n_100),
	.Q(n_406),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44816 (.A(DPATH_RF_MEMORY_7__29_),
	.B(n_98),
	.Q(n_405),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44817 (.A(DPATH_RF_MEMORY_7__30_),
	.B(n_96),
	.Q(n_404),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44818 (.A(DPATH_RF_MEMORY_7__31_),
	.B(n_94),
	.Q(n_403),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g44819 (.A(DPATH_RF_MEMORY_1__3_),
	.B(n_143),
	.Q(n_402),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44820 (.A(DPATH_RF_MEMORY_9__1_),
	.B(n_139),
	.Q(n_401),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44821 (.A(DPATH_RF_MEMORY_9__0_),
	.B(n_116),
	.Q(n_400),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44822 (.A(DPATH_RF_MEMORY_9__3_),
	.B(n_143),
	.Q(n_399),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44823 (.A(DPATH_RF_MEMORY_9__5_),
	.B(n_151),
	.Q(n_398),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44824 (.A(DPATH_RF_MEMORY_9__7_),
	.B(n_106),
	.Q(n_397),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44825 (.A(DPATH_RF_MEMORY_9__8_),
	.B(n_135),
	.Q(n_396),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44826 (.A(DPATH_RF_MEMORY_9__9_),
	.B(n_120),
	.Q(n_395),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44827 (.A(DPATH_RF_MEMORY_9__11_),
	.B(n_131),
	.Q(n_394),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44828 (.A(DPATH_RF_MEMORY_9__12_),
	.B(n_129),
	.Q(n_393),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44829 (.A(DPATH_RF_MEMORY_9__13_),
	.B(n_141),
	.Q(n_392),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44830 (.A(DPATH_RF_MEMORY_9__14_),
	.B(n_126),
	.Q(n_391),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44831 (.A(DPATH_RF_MEMORY_9__16_),
	.B(n_153),
	.Q(n_390),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44832 (.A(DPATH_RF_MEMORY_1__0_),
	.B(n_116),
	.Q(n_389),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44833 (.A(DPATH_RF_MEMORY_9__17_),
	.B(n_118),
	.Q(n_388),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44834 (.A(DPATH_RF_MEMORY_9__15_),
	.B(n_124),
	.Q(n_387),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44835 (.A(DPATH_RF_MEMORY_9__18_),
	.B(n_147),
	.Q(n_386),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44836 (.A(DPATH_RF_MEMORY_9__19_),
	.B(n_114),
	.Q(n_385),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44837 (.A(DPATH_RF_MEMORY_9__20_),
	.B(n_112),
	.Q(n_384),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44838 (.A(DPATH_RF_MEMORY_9__21_),
	.B(n_145),
	.Q(n_383),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44839 (.A(DPATH_RF_MEMORY_9__22_),
	.B(n_149),
	.Q(n_382),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44840 (.A(DPATH_RF_MEMORY_9__23_),
	.B(n_122),
	.Q(n_381),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44841 (.A(DPATH_RF_MEMORY_9__24_),
	.B(n_110),
	.Q(n_380),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44842 (.A(DPATH_RF_MEMORY_9__25_),
	.B(n_108),
	.Q(n_379),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44843 (.A(DPATH_RF_MEMORY_9__26_),
	.B(n_104),
	.Q(n_378),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44844 (.A(DPATH_RF_MEMORY_9__27_),
	.B(n_102),
	.Q(n_377),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44845 (.A(DPATH_RF_MEMORY_9__28_),
	.B(n_100),
	.Q(n_376),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44846 (.A(DPATH_RF_MEMORY_9__29_),
	.B(n_98),
	.Q(n_375),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44847 (.A(DPATH_RF_MEMORY_1__1_),
	.B(n_139),
	.Q(n_374),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44848 (.A(DPATH_RF_MEMORY_9__31_),
	.B(n_94),
	.Q(n_373),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44849 (.A(DPATH_RF_MEMORY_1__4_),
	.B(n_92),
	.Q(n_372),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44850 (.A(DPATH_RF_MEMORY_1__5_),
	.B(n_151),
	.Q(n_371),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44851 (.A(DPATH_RF_MEMORY_9__30_),
	.B(n_96),
	.Q(n_370),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44852 (.A(DPATH_RF_MEMORY_1__6_),
	.B(n_137),
	.Q(n_369),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44853 (.A(DPATH_RF_MEMORY_1__7_),
	.B(n_106),
	.Q(n_368),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44854 (.A(DPATH_RF_MEMORY_1__8_),
	.B(n_135),
	.Q(n_367),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44855 (.A(DPATH_RF_MEMORY_11__0_),
	.B(n_116),
	.Q(n_366),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44856 (.A(DPATH_RF_MEMORY_11__1_),
	.B(n_139),
	.Q(n_365),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44857 (.A(DPATH_RF_MEMORY_1__9_),
	.B(n_120),
	.Q(n_364),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44858 (.A(DPATH_RF_MEMORY_11__3_),
	.B(n_143),
	.Q(n_363),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44859 (.A(DPATH_RF_MEMORY_11__4_),
	.B(n_92),
	.Q(n_362),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44860 (.A(DPATH_RF_MEMORY_11__5_),
	.B(n_151),
	.Q(n_361),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44861 (.A(DPATH_RF_MEMORY_11__6_),
	.B(n_137),
	.Q(n_360),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44862 (.A(DPATH_RF_MEMORY_11__7_),
	.B(n_106),
	.Q(n_359),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44863 (.A(DPATH_RF_MEMORY_11__8_),
	.B(n_135),
	.Q(n_358),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44864 (.A(DPATH_RF_MEMORY_11__9_),
	.B(n_120),
	.Q(n_357),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44865 (.A(DPATH_RF_MEMORY_1__11_),
	.B(n_131),
	.Q(n_356),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44866 (.A(DPATH_RF_MEMORY_11__10_),
	.B(n_133),
	.Q(n_355),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44867 (.A(DPATH_RF_MEMORY_1__10_),
	.B(n_133),
	.Q(n_354),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44868 (.A(DPATH_RF_MEMORY_11__11_),
	.B(n_131),
	.Q(n_353),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44869 (.A(DPATH_RF_MEMORY_11__12_),
	.B(n_129),
	.Q(n_352),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44870 (.A(DPATH_RF_MEMORY_11__13_),
	.B(n_141),
	.Q(n_351),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44871 (.A(DPATH_RF_MEMORY_1__13_),
	.B(n_141),
	.Q(n_350),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44872 (.A(DPATH_RF_MEMORY_11__14_),
	.B(n_126),
	.Q(n_349),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44873 (.A(DPATH_RF_MEMORY_11__15_),
	.B(n_124),
	.Q(n_348),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44874 (.A(DPATH_RF_MEMORY_11__16_),
	.B(n_153),
	.Q(n_347),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44875 (.A(DPATH_RF_MEMORY_11__17_),
	.B(n_118),
	.Q(n_346),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44876 (.A(DPATH_RF_MEMORY_11__18_),
	.B(n_147),
	.Q(n_345),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44877 (.A(DPATH_RF_MEMORY_11__19_),
	.B(n_114),
	.Q(n_344),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44878 (.A(DPATH_RF_MEMORY_11__20_),
	.B(n_112),
	.Q(n_343),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44879 (.A(DPATH_RF_MEMORY_11__21_),
	.B(n_145),
	.Q(n_342),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44880 (.A(DPATH_RF_MEMORY_11__22_),
	.B(n_149),
	.Q(n_341),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44881 (.A(DPATH_RF_MEMORY_1__14_),
	.B(n_126),
	.Q(n_340),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44882 (.A(DPATH_RF_MEMORY_11__23_),
	.B(n_122),
	.Q(n_339),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44883 (.A(DPATH_RF_MEMORY_11__24_),
	.B(n_110),
	.Q(n_338),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44884 (.A(DPATH_RF_MEMORY_11__25_),
	.B(n_108),
	.Q(n_337),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44885 (.A(DPATH_RF_MEMORY_11__26_),
	.B(n_104),
	.Q(n_336),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44886 (.A(DPATH_RF_MEMORY_1__12_),
	.B(n_129),
	.Q(n_335),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44887 (.A(DPATH_RF_MEMORY_11__27_),
	.B(n_102),
	.Q(n_334),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44888 (.A(DPATH_RF_MEMORY_1__15_),
	.B(n_124),
	.Q(n_333),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44889 (.A(DPATH_RF_MEMORY_11__28_),
	.B(n_100),
	.Q(n_332),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44890 (.A(DPATH_RF_MEMORY_11__29_),
	.B(n_98),
	.Q(n_331),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44891 (.A(DPATH_RF_MEMORY_11__30_),
	.B(n_96),
	.Q(n_330),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44892 (.A(DPATH_RF_MEMORY_11__31_),
	.B(n_94),
	.Q(n_329),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g44893 (.A(DPATH_RF_MEMORY_1__16_),
	.B(n_153),
	.Q(n_328),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44894 (.A(DPATH_RF_MEMORY_1__17_),
	.B(n_118),
	.Q(n_327),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44895 (.A(DPATH_RF_MEMORY_1__18_),
	.B(n_147),
	.Q(n_326),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44896 (.A(DPATH_RF_MEMORY_1__19_),
	.B(n_114),
	.Q(n_325),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44897 (.A(DPATH_RF_MEMORY_1__20_),
	.B(n_112),
	.Q(n_324),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44898 (.A(DPATH_RF_MEMORY_1__21_),
	.B(n_145),
	.Q(n_323),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44899 (.A(DPATH_RF_MEMORY_1__22_),
	.B(n_149),
	.Q(n_322),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44900 (.A(DPATH_RF_MEMORY_1__23_),
	.B(n_122),
	.Q(n_321),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44901 (.A(DPATH_RF_MEMORY_1__24_),
	.B(n_110),
	.Q(n_320),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44902 (.A(DPATH_RF_MEMORY_1__25_),
	.B(n_108),
	.Q(n_319),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44903 (.A(DPATH_RF_MEMORY_1__27_),
	.B(n_102),
	.Q(n_318),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44904 (.A(DPATH_RF_MEMORY_1__28_),
	.B(n_100),
	.Q(n_317),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44905 (.A(DPATH_RF_MEMORY_1__29_),
	.B(n_98),
	.Q(n_316),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44906 (.A(DPATH_RF_MEMORY_1__26_),
	.B(n_104),
	.Q(n_315),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44907 (.A(DPATH_RF_MEMORY_1__30_),
	.B(n_96),
	.Q(n_314),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44908 (.A(DPATH_RF_MEMORY_1__31_),
	.B(n_94),
	.Q(n_313),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g44909 (.A(DPATH_RF_MEMORY_15__0_),
	.B(n_116),
	.Q(n_312),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44910 (.A(DPATH_RF_MEMORY_15__1_),
	.B(n_139),
	.Q(n_311),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44911 (.A(DPATH_RF_MEMORY_15__3_),
	.B(n_143),
	.Q(n_310),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44912 (.A(DPATH_RF_MEMORY_15__4_),
	.B(n_92),
	.Q(n_309),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44913 (.A(DPATH_RF_MEMORY_15__5_),
	.B(n_151),
	.Q(n_308),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44914 (.A(DPATH_RF_MEMORY_15__6_),
	.B(n_137),
	.Q(n_307),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44915 (.A(DPATH_RF_MEMORY_15__7_),
	.B(n_106),
	.Q(n_306),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44916 (.A(DPATH_RF_MEMORY_15__8_),
	.B(n_135),
	.Q(n_305),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44917 (.A(DPATH_RF_MEMORY_15__9_),
	.B(n_120),
	.Q(n_304),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44918 (.A(DPATH_RF_MEMORY_15__10_),
	.B(n_133),
	.Q(n_303),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44919 (.A(DPATH_RF_MEMORY_15__11_),
	.B(n_131),
	.Q(n_302),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44920 (.A(DPATH_RF_MEMORY_15__12_),
	.B(n_129),
	.Q(n_301),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44921 (.A(DPATH_RF_MEMORY_15__13_),
	.B(n_141),
	.Q(n_300),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44922 (.A(DPATH_RF_MEMORY_15__14_),
	.B(n_126),
	.Q(n_299),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44923 (.A(DPATH_RF_MEMORY_15__15_),
	.B(n_124),
	.Q(n_298),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44924 (.A(DPATH_RF_MEMORY_15__16_),
	.B(n_153),
	.Q(n_297),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44925 (.A(DPATH_RF_MEMORY_15__17_),
	.B(n_118),
	.Q(n_296),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44926 (.A(DPATH_RF_MEMORY_15__18_),
	.B(n_147),
	.Q(n_295),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44927 (.A(DPATH_RF_MEMORY_15__19_),
	.B(n_114),
	.Q(n_294),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44928 (.A(DPATH_RF_MEMORY_15__20_),
	.B(n_112),
	.Q(n_293),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44929 (.A(DPATH_RF_MEMORY_15__21_),
	.B(n_145),
	.Q(n_292),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44930 (.A(DPATH_RF_MEMORY_15__22_),
	.B(n_149),
	.Q(n_291),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44931 (.A(DPATH_RF_MEMORY_15__23_),
	.B(n_122),
	.Q(n_290),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44932 (.A(DPATH_RF_MEMORY_15__24_),
	.B(n_110),
	.Q(n_289),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44933 (.A(DPATH_RF_MEMORY_15__25_),
	.B(n_108),
	.Q(n_288),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44934 (.A(DPATH_RF_MEMORY_15__26_),
	.B(n_104),
	.Q(n_287),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44935 (.A(DPATH_RF_MEMORY_15__27_),
	.B(n_102),
	.Q(n_286),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44936 (.A(DPATH_RF_MEMORY_15__28_),
	.B(n_100),
	.Q(n_285),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44937 (.A(DPATH_RF_MEMORY_15__29_),
	.B(n_98),
	.Q(n_284),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44938 (.A(DPATH_RF_MEMORY_9__10_),
	.B(n_133),
	.Q(n_283),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44939 (.A(DPATH_RF_MEMORY_15__30_),
	.B(n_96),
	.Q(n_282),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44940 (.A(DPATH_RF_MEMORY_15__31_),
	.B(n_94),
	.Q(n_281),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g44941 (.A(DPATH_RF_MEMORY_3__0_),
	.B(n_116),
	.Q(n_280),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44942 (.A(DPATH_RF_MEMORY_3__1_),
	.B(n_139),
	.Q(n_279),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44943 (.A(DPATH_RF_MEMORY_3__4_),
	.B(n_92),
	.Q(n_278),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44944 (.A(DPATH_RF_MEMORY_3__3_),
	.B(n_143),
	.Q(n_277),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44945 (.A(DPATH_RF_MEMORY_3__5_),
	.B(n_151),
	.Q(n_276),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44946 (.A(DPATH_RF_MEMORY_3__6_),
	.B(n_137),
	.Q(n_275),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44947 (.A(DPATH_RF_MEMORY_3__7_),
	.B(n_106),
	.Q(n_274),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44948 (.A(DPATH_RF_MEMORY_3__8_),
	.B(n_135),
	.Q(n_273),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44949 (.A(DPATH_RF_MEMORY_3__9_),
	.B(n_120),
	.Q(n_272),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44950 (.A(DPATH_RF_MEMORY_3__10_),
	.B(n_133),
	.Q(n_271),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44951 (.A(DPATH_RF_MEMORY_3__11_),
	.B(n_131),
	.Q(n_270),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44952 (.A(DPATH_RF_MEMORY_17__0_),
	.B(n_116),
	.Q(n_269),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44953 (.A(DPATH_RF_MEMORY_3__12_),
	.B(n_129),
	.Q(n_268),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44954 (.A(DPATH_RF_MEMORY_17__1_),
	.B(n_139),
	.Q(n_267),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44955 (.A(DPATH_RF_MEMORY_3__13_),
	.B(n_141),
	.Q(n_266),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44956 (.A(DPATH_RF_MEMORY_17__3_),
	.B(n_143),
	.Q(n_265),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44957 (.A(DPATH_RF_MEMORY_17__4_),
	.B(n_92),
	.Q(n_264),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44958 (.A(DPATH_RF_MEMORY_17__5_),
	.B(n_151),
	.Q(n_263),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44959 (.A(DPATH_RF_MEMORY_3__14_),
	.B(n_126),
	.Q(n_262),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44960 (.A(DPATH_RF_MEMORY_17__6_),
	.B(n_137),
	.Q(n_261),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44961 (.A(DPATH_RF_MEMORY_3__15_),
	.B(n_124),
	.Q(n_260),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44962 (.A(DPATH_RF_MEMORY_17__7_),
	.B(n_106),
	.Q(n_259),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44963 (.A(DPATH_RF_MEMORY_9__6_),
	.B(n_137),
	.Q(n_258),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44964 (.A(DPATH_RF_MEMORY_3__16_),
	.B(n_153),
	.Q(n_257),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44965 (.A(DPATH_RF_MEMORY_17__8_),
	.B(n_135),
	.Q(n_256),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44966 (.A(DPATH_RF_MEMORY_17__9_),
	.B(n_120),
	.Q(n_255),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44967 (.A(DPATH_RF_MEMORY_17__10_),
	.B(n_133),
	.Q(n_254),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44968 (.A(DPATH_RF_MEMORY_3__17_),
	.B(n_118),
	.Q(n_253),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44969 (.A(DPATH_RF_MEMORY_17__11_),
	.B(n_131),
	.Q(n_252),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44970 (.A(DPATH_RF_MEMORY_3__18_),
	.B(n_147),
	.Q(n_251),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44971 (.A(DPATH_RF_MEMORY_17__12_),
	.B(n_129),
	.Q(n_250),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44972 (.A(DPATH_RF_MEMORY_17__13_),
	.B(n_141),
	.Q(n_249),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44973 (.A(DPATH_RF_MEMORY_17__14_),
	.B(n_126),
	.Q(n_248),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44974 (.A(DPATH_RF_MEMORY_17__15_),
	.B(n_124),
	.Q(n_247),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44975 (.A(DPATH_RF_MEMORY_9__4_),
	.B(n_92),
	.Q(n_246),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g44976 (.A(DPATH_RF_MEMORY_17__16_),
	.B(n_153),
	.Q(n_245),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44977 (.A(DPATH_RF_MEMORY_3__19_),
	.B(n_114),
	.Q(n_244),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44978 (.A(DPATH_RF_MEMORY_17__17_),
	.B(n_118),
	.Q(n_243),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44979 (.A(DPATH_RF_MEMORY_3__20_),
	.B(n_112),
	.Q(n_242),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44980 (.A(DPATH_RF_MEMORY_17__18_),
	.B(n_147),
	.Q(n_241),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44981 (.A(DPATH_RF_MEMORY_3__21_),
	.B(n_145),
	.Q(n_240),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44982 (.A(DPATH_RF_MEMORY_17__19_),
	.B(n_114),
	.Q(n_239),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44983 (.A(DPATH_RF_MEMORY_17__20_),
	.B(n_112),
	.Q(n_238),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44984 (.A(DPATH_RF_MEMORY_17__21_),
	.B(n_145),
	.Q(n_237),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44985 (.A(DPATH_RF_MEMORY_3__22_),
	.B(n_149),
	.Q(n_236),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44986 (.A(DPATH_RF_MEMORY_17__22_),
	.B(n_149),
	.Q(n_235),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44987 (.A(DPATH_RF_MEMORY_3__23_),
	.B(n_122),
	.Q(n_234),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44988 (.A(DPATH_RF_MEMORY_17__23_),
	.B(n_122),
	.Q(n_233),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44989 (.A(DPATH_RF_MEMORY_3__24_),
	.B(n_110),
	.Q(n_232),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44990 (.A(DPATH_RF_MEMORY_17__24_),
	.B(n_110),
	.Q(n_231),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44991 (.A(DPATH_RF_MEMORY_17__25_),
	.B(n_108),
	.Q(n_230),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44992 (.A(DPATH_RF_MEMORY_17__26_),
	.B(n_104),
	.Q(n_229),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44993 (.A(DPATH_RF_MEMORY_3__25_),
	.B(n_108),
	.Q(n_228),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44994 (.A(DPATH_RF_MEMORY_17__27_),
	.B(n_102),
	.Q(n_227),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44995 (.A(DPATH_RF_MEMORY_17__28_),
	.B(n_100),
	.Q(n_226),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44996 (.A(DPATH_RF_MEMORY_3__26_),
	.B(n_104),
	.Q(n_225),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44997 (.A(DPATH_RF_MEMORY_17__29_),
	.B(n_98),
	.Q(n_224),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g44998 (.A(DPATH_RF_MEMORY_3__27_),
	.B(n_102),
	.Q(n_223),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g44999 (.A(DPATH_RF_MEMORY_17__30_),
	.B(n_96),
	.Q(n_222),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g45000 (.A(DPATH_RF_MEMORY_17__31_),
	.B(n_94),
	.Q(n_221),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g45001 (.A(DPATH_RF_MEMORY_3__28_),
	.B(n_100),
	.Q(n_220),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g45002 (.A(DPATH_RF_MEMORY_3__29_),
	.B(n_98),
	.Q(n_219),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g45003 (.A(DPATH_RF_MEMORY_3__30_),
	.B(n_96),
	.Q(n_218),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g45004 (.A(DPATH_RF_MEMORY_3__31_),
	.B(n_94),
	.Q(n_217),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g45005 (.A(DPATH_RF_MEMORY_19__0_),
	.B(n_116),
	.Q(n_216),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45006 (.A(DPATH_RF_MEMORY_19__1_),
	.B(n_139),
	.Q(n_215),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45007 (.A(DPATH_RF_MEMORY_19__3_),
	.B(n_143),
	.Q(n_214),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45008 (.A(DPATH_RF_MEMORY_19__4_),
	.B(n_92),
	.Q(n_213),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45009 (.A(DPATH_RF_MEMORY_19__5_),
	.B(n_151),
	.Q(n_212),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45010 (.A(DPATH_RF_MEMORY_19__6_),
	.B(n_137),
	.Q(n_211),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45011 (.A(DPATH_RF_MEMORY_19__7_),
	.B(n_106),
	.Q(n_210),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45012 (.A(DPATH_RF_MEMORY_19__8_),
	.B(n_135),
	.Q(n_209),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45013 (.A(DPATH_RF_MEMORY_19__9_),
	.B(n_120),
	.Q(n_208),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45014 (.A(DPATH_RF_MEMORY_19__10_),
	.B(n_133),
	.Q(n_207),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45015 (.A(DPATH_RF_MEMORY_19__11_),
	.B(n_131),
	.Q(n_206),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45016 (.A(DPATH_RF_MEMORY_19__12_),
	.B(n_129),
	.Q(n_205),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45017 (.A(DPATH_RF_MEMORY_19__13_),
	.B(n_141),
	.Q(n_204),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45018 (.A(DPATH_RF_MEMORY_19__14_),
	.B(n_126),
	.Q(n_203),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45019 (.A(DPATH_RF_MEMORY_19__15_),
	.B(n_124),
	.Q(n_202),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45020 (.A(DPATH_RF_MEMORY_19__16_),
	.B(n_153),
	.Q(n_201),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45021 (.A(DPATH_RF_MEMORY_19__17_),
	.B(n_118),
	.Q(n_200),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45022 (.A(DPATH_RF_MEMORY_19__18_),
	.B(n_147),
	.Q(n_199),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45023 (.A(DPATH_RF_MEMORY_19__19_),
	.B(n_114),
	.Q(n_198),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45024 (.A(DPATH_RF_MEMORY_19__20_),
	.B(n_112),
	.Q(n_197),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45025 (.A(DPATH_RF_MEMORY_19__21_),
	.B(n_145),
	.Q(n_196),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45026 (.A(DPATH_RF_MEMORY_19__22_),
	.B(n_149),
	.Q(n_195),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45027 (.A(DPATH_RF_MEMORY_19__23_),
	.B(n_122),
	.Q(n_194),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45028 (.A(DPATH_RF_MEMORY_19__24_),
	.B(n_110),
	.Q(n_193),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45029 (.A(DPATH_RF_MEMORY_19__25_),
	.B(n_108),
	.Q(n_192),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45030 (.A(DPATH_RF_MEMORY_19__26_),
	.B(n_104),
	.Q(n_191),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45031 (.A(DPATH_RF_MEMORY_19__27_),
	.B(n_102),
	.Q(n_190),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45032 (.A(DPATH_RF_MEMORY_19__28_),
	.B(n_100),
	.Q(n_189),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45033 (.A(DPATH_RF_MEMORY_19__29_),
	.B(n_98),
	.Q(n_188),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45034 (.A(DPATH_RF_MEMORY_19__30_),
	.B(n_96),
	.Q(n_187),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45035 (.A(DPATH_RF_MEMORY_19__31_),
	.B(n_94),
	.Q(n_186),
	.S0(FE_OFN21_n_89));
   MUX2_X2_50_SVT g45036 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_22__2_),
	.Q(n_185),
	.S0(n_72));
   MUX2_X2_50_SVT g45037 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_24__2_),
	.Q(n_184),
	.S0(n_86));
   MUX2_X2_50_SVT g45038 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_25__2_),
	.Q(n_183),
	.S0(FE_OFN0_n_2));
   MUX2_X2_50_SVT g45039 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_26__2_),
	.Q(n_182),
	.S0(n_82));
   MUX2_X2_50_SVT g45040 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_8__2_),
	.Q(n_181),
	.S0(FE_OFN15_n_83));
   MUX2_X2_50_SVT g45041 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_28__2_),
	.Q(n_180),
	.S0(n_85));
   MUX2_X2_50_SVT g45042 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_29__2_),
	.Q(n_179),
	.S0(n_67));
   MUX2_X2_50_SVT g45043 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_30__2_),
	.Q(n_178),
	.S0(FE_OFN78_n_79));
   MUX2_X2_50_SVT g45044 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_10__2_),
	.Q(n_177),
	.S0(n_81));
   MUX2_X2_50_SVT g45045 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_12__2_),
	.Q(n_176),
	.S0(n_62));
   MUX2_X2_50_SVT g45046 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_14__2_),
	.Q(n_175),
	.S0(FE_OFN5_n_69));
   MUX2_X2_50_SVT g45047 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_16__2_),
	.Q(n_174),
	.S0(FE_OFN75_n_73));
   MUX2_X2_50_SVT g45048 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_18__2_),
	.Q(n_173),
	.S0(FE_OFN76_n_75));
   MUX2_X2_50_SVT g45049 (.A(FE_OFN101_n_128),
	.B(DPATH_RF_MEMORY_4__2_),
	.Q(n_172),
	.S0(FE_OFN3_n_64));
   MUX2_X2_50_SVT g45050 (.A(n_128),
	.B(DPATH_RF_MEMORY_20__2_),
	.Q(n_171),
	.S0(n_76));
   MUX2_X2_50_SVT g45051 (.A(DPATH_RF_MEMORY_6__2_),
	.B(FE_OFN101_n_128),
	.Q(n_170),
	.S0(n_65));
   MUX2_X2_50_SVT g45052 (.A(DPATH_RF_MEMORY_27__2_),
	.B(FE_OFN101_n_128),
	.Q(n_169),
	.S0(n_66));
   MUX2_X2_50_SVT g45053 (.A(DPATH_RF_MEMORY_31__2_),
	.B(FE_OFN101_n_128),
	.Q(n_168),
	.S0(n_68));
   MUX2_X2_50_SVT g45054 (.A(DPATH_RF_MEMORY_2__2_),
	.B(FE_OFN101_n_128),
	.Q(n_167),
	.S0(n_63));
   MUX2_X2_50_SVT g45055 (.A(DPATH_RF_MEMORY_13__2_),
	.B(FE_OFN101_n_128),
	.Q(n_166),
	.S0(FE_OFN23_n_91));
   MUX2_X2_50_SVT g45056 (.A(DPATH_RF_MEMORY_5__2_),
	.B(FE_OFN101_n_128),
	.Q(n_165),
	.S0(FE_OFN9_n_74));
   MUX2_X2_50_SVT g45057 (.A(DPATH_RF_MEMORY_21__2_),
	.B(FE_OFN101_n_128),
	.Q(n_164),
	.S0(FE_OFN13_n_80));
   MUX2_X2_50_SVT g45058 (.A(DPATH_RF_MEMORY_23__2_),
	.B(FE_OFN101_n_128),
	.Q(n_163),
	.S0(FE_OFN16_n_84));
   MUX2_X2_50_SVT g45059 (.A(DPATH_RF_MEMORY_7__2_),
	.B(FE_OFN101_n_128),
	.Q(n_162),
	.S0(FE_OFN17_n_87));
   MUX2_X2_50_SVT g45060 (.A(DPATH_RF_MEMORY_1__2_),
	.B(FE_OFN101_n_128),
	.Q(n_161),
	.S0(FE_OFN10_n_77));
   MUX2_X2_50_SVT g45061 (.A(DPATH_RF_MEMORY_11__2_),
	.B(FE_OFN101_n_128),
	.Q(n_160),
	.S0(FE_OFN12_n_78));
   MUX2_X2_50_SVT g45062 (.A(DPATH_RF_MEMORY_15__2_),
	.B(FE_OFN101_n_128),
	.Q(n_159),
	.S0(FE_OFN22_n_90));
   MUX2_X2_50_SVT g45063 (.A(DPATH_RF_MEMORY_3__2_),
	.B(FE_OFN101_n_128),
	.Q(n_158),
	.S0(FE_OFN19_n_88));
   MUX2_X2_50_SVT g45064 (.A(DPATH_RF_MEMORY_17__2_),
	.B(n_128),
	.Q(n_157),
	.S0(FE_OFN6_n_70));
   MUX2_X2_50_SVT g45065 (.A(DPATH_RF_MEMORY_9__2_),
	.B(FE_OFN101_n_128),
	.Q(n_156),
	.S0(FE_OFN8_n_71));
   MUX2_X2_50_SVT g45066 (.A(DPATH_RF_MEMORY_19__2_),
	.B(n_128),
	.Q(n_155),
	.S0(FE_OFN21_n_89));
   INV_X2_50_SVT g45099 (.A(FE_OFN117_n_154),
	.Q(n_153));
   INV_X2_50_SVT g45100 (.A(FE_OFN116_n_152),
	.Q(n_151));
   INV_X2_50_SVT g45101 (.A(FE_OFN114_n_150),
	.Q(n_149));
   INV_X2_50_SVT g45103 (.A(FE_OFN112_n_146),
	.Q(n_145));
   INV_X2_50_SVT g45104 (.A(FE_OFN111_n_144),
	.Q(n_143));
   INV_X2_50_SVT g45105 (.A(FE_OFN110_n_142),
	.Q(n_141));
   INV_X2_50_SVT g45107 (.A(FE_OFN107_n_138),
	.Q(n_137));
   INV_X2_50_SVT g45108 (.A(FE_OFN106_n_136),
	.Q(n_135));
   INV_X2_50_SVT g45109 (.A(FE_OFN105_n_134),
	.Q(n_133));
   INV_X2_50_SVT g45111 (.A(FE_OFN102_n_130),
	.Q(n_129));
   INV_X2_50_SVT g45112 (.A(FE_OFN100_n_127),
	.Q(n_126));
   INV_X2_50_SVT g45113 (.A(FE_OFN99_n_125),
	.Q(n_124));
   INV_X2_50_SVT g45114 (.A(FE_OFN97_n_123),
	.Q(n_122));
   INV_X2_50_SVT g45115 (.A(FE_OFN96_n_121),
	.Q(n_120));
   INV_X2_50_SVT g45116 (.A(FE_OFN95_n_119),
	.Q(n_118));
   INV_X2_50_SVT g45117 (.A(FE_OFN93_n_117),
	.Q(n_116));
   INV_X2_50_SVT g45120 (.A(FE_OFN90_n_111),
	.Q(n_110));
   INV_X2_50_SVT g45122 (.A(FE_OFN88_n_107),
	.Q(n_106));
   INV_X2_50_SVT g45123 (.A(FE_OFN87_n_105),
	.Q(n_104));
   INV_X2_50_SVT g45126 (.A(FE_OFN84_n_99),
	.Q(n_98));
   INV_X2_50_SVT g45127 (.A(FE_OFN83_n_97),
	.Q(n_96));
   AOI222_X0_50_SVT g45130 (.A0(ALURSLT[16]),
	.A1(n_0),
	.B0(DPATH_n_2876),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[16]),
	.Q(n_154));
   AOI222_X0_50_SVT g45131 (.A0(ALURSLT[5]),
	.A1(n_0),
	.B0(DPATH_n_2887),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[5]),
	.Q(n_152));
   AOI222_X0_50_SVT g45132 (.A0(ALURSLT[22]),
	.A1(n_0),
	.B0(DPATH_n_2870),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[22]),
	.Q(n_150));
   AOI222_X0_50_SVT g45133 (.A0(ALURSLT[18]),
	.A1(n_0),
	.B0(DPATH_n_2874),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[18]),
	.Q(n_148));
   AOI222_X0_50_SVT g45134 (.A0(ALURSLT[21]),
	.A1(n_0),
	.B0(DPATH_n_2871),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[21]),
	.Q(n_146));
   AOI222_X0_50_SVT g45135 (.A0(ALURSLT[3]),
	.A1(n_0),
	.B0(DPATH_n_2889),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[3]),
	.Q(n_144));
   AOI222_X0_50_SVT g45136 (.A0(ALURSLT[13]),
	.A1(n_0),
	.B0(DPATH_n_2879),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[13]),
	.Q(n_142));
   AOI222_X0_50_SVT g45137 (.A0(ALURSLT[1]),
	.A1(n_0),
	.B0(PC[1]),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[1]),
	.Q(n_140));
   AOI222_X0_50_SVT g45138 (.A0(ALURSLT[6]),
	.A1(n_0),
	.B0(DPATH_n_2886),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[6]),
	.Q(n_138));
   AOI222_X0_50_SVT g45139 (.A0(ALURSLT[8]),
	.A1(n_0),
	.B0(DPATH_n_2884),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[8]),
	.Q(n_136));
   AOI222_X0_50_SVT g45140 (.A0(ALURSLT[10]),
	.A1(n_0),
	.B0(DPATH_n_2882),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[10]),
	.Q(n_134));
   AOI222_X0_50_SVT g45141 (.A0(ALURSLT[11]),
	.A1(n_0),
	.B0(DPATH_n_2881),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[11]),
	.Q(n_132));
   AOI222_X0_50_SVT g45142 (.A0(ALURSLT[12]),
	.A1(n_0),
	.B0(DPATH_n_2880),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[12]),
	.Q(n_130));
   NAND2_A_NAND2_X1_50_SVT g45143 (.A0N(n_4),
	.A1N(DMEMRD[2]),
	.B0(n_61),
	.Q(n_128));
   AOI222_X0_50_SVT g45144 (.A0(ALURSLT[14]),
	.A1(n_0),
	.B0(DPATH_n_2878),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[14]),
	.Q(n_127));
   AOI222_X0_50_SVT g45145 (.A0(ALURSLT[15]),
	.A1(n_0),
	.B0(DPATH_n_2877),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[15]),
	.Q(n_125));
   AOI222_X0_50_SVT g45146 (.A0(ALURSLT[23]),
	.A1(n_0),
	.B0(DPATH_n_2869),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[23]),
	.Q(n_123));
   AOI222_X0_50_SVT g45147 (.A0(ALURSLT[9]),
	.A1(n_0),
	.B0(DPATH_n_2883),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[9]),
	.Q(n_121));
   AOI222_X0_50_SVT g45148 (.A0(ALURSLT[17]),
	.A1(n_0),
	.B0(DPATH_n_2875),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[17]),
	.Q(n_119));
   AOI222_X0_50_SVT g45149 (.A0(ALURSLT[0]),
	.A1(n_0),
	.B0(PC[0]),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[0]),
	.Q(n_117));
   AOI222_X0_50_SVT g45150 (.A0(ALURSLT[19]),
	.A1(n_0),
	.B0(DPATH_n_2873),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[19]),
	.Q(n_115));
   AOI222_X0_50_SVT g45151 (.A0(ALURSLT[20]),
	.A1(n_0),
	.B0(DPATH_n_2872),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[20]),
	.Q(n_113));
   AOI222_X0_50_SVT g45152 (.A0(ALURSLT[24]),
	.A1(n_0),
	.B0(DPATH_n_2868),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[24]),
	.Q(n_111));
   AOI222_X0_50_SVT g45153 (.A0(ALURSLT[25]),
	.A1(n_0),
	.B0(DPATH_n_2867),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[25]),
	.Q(n_109));
   AOI222_X0_50_SVT g45154 (.A0(ALURSLT[7]),
	.A1(n_0),
	.B0(DPATH_n_2885),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[7]),
	.Q(n_107));
   AOI222_X0_50_SVT g45155 (.A0(ALURSLT[26]),
	.A1(n_0),
	.B0(DPATH_n_2866),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[26]),
	.Q(n_105));
   AOI222_X0_50_SVT g45156 (.A0(ALURSLT[27]),
	.A1(n_0),
	.B0(DPATH_n_2865),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[27]),
	.Q(n_103));
   AOI222_X0_50_SVT g45157 (.A0(ALURSLT[28]),
	.A1(n_0),
	.B0(DPATH_n_2864),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[28]),
	.Q(n_101));
   AOI222_X0_50_SVT g45158 (.A0(ALURSLT[29]),
	.A1(n_0),
	.B0(DPATH_n_2863),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[29]),
	.Q(n_99));
   AOI222_X0_50_SVT g45159 (.A0(ALURSLT[30]),
	.A1(n_0),
	.B0(DPATH_n_2862),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[30]),
	.Q(n_97));
   AOI222_X0_50_SVT g45160 (.A0(ALURSLT[31]),
	.A1(n_0),
	.B0(DPATH_n_2861),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[31]),
	.Q(n_95));
   AOI222_X0_50_SVT g45161 (.A0(ALURSLT[4]),
	.A1(n_0),
	.B0(DPATH_n_2888),
	.B1(INSTR[2]),
	.C0(n_4),
	.C1(DMEMRD[4]),
	.Q(n_93));
   NOR2_A_AOI21_X2_50_SVT g45162 (.A0N(PC[2]),
	.A1N(n_3),
	.B0(ALURSLT[2]),
	.B1(n_0),
	.Q(n_61));
   NOR2_X0_50_SVT g45163 (.A(n_22),
	.B(n_14),
	.Q(n_91));
   NOR2_X0_50_SVT g45164 (.A(n_26),
	.B(n_14),
	.Q(n_90));
   NOR2_X0_50_SVT g45165 (.A(n_24),
	.B(n_13),
	.Q(n_89));
   NOR2_X0_50_SVT g45166 (.A(n_24),
	.B(n_16),
	.Q(n_88));
   NOR2_X0_50_SVT g45167 (.A(n_26),
	.B(n_16),
	.Q(n_87));
   NAND2_X1_50_SVT g45168 (.A(n_27),
	.B(n_17),
	.Q(n_86));
   NAND2_X2_50_SVT g45169 (.A(n_21),
	.B(n_17),
	.Q(n_85));
   NOR2_X0_50_SVT g45170 (.A(n_26),
	.B(n_13),
	.Q(n_84));
   NAND2_X0_50_SVT g45171 (.A(n_27),
	.B(n_1),
	.Q(n_83));
   CLKNAND2_X4_50_SVT g45172 (.A(n_23),
	.B(n_17),
	.Q(n_82));
   NAND2_X6_50_SVT g45173 (.A(n_23),
	.B(n_1),
	.Q(n_81));
   NOR2_X0_50_SVT g45174 (.A(n_22),
	.B(n_13),
	.Q(n_80));
   NAND2_X0_50_SVT g45175 (.A(n_25),
	.B(n_17),
	.Q(n_79));
   NOR2_X0_50_SVT g45176 (.A(n_24),
	.B(n_14),
	.Q(n_78));
   NOR2_X0_50_SVT g45177 (.A(n_28),
	.B(n_16),
	.Q(n_77));
   CLKNAND2_X2_50_SVT g45178 (.A(n_21),
	.B(n_15),
	.Q(n_76));
   NAND2_X0_50_SVT g45179 (.A(n_23),
	.B(n_15),
	.Q(n_75));
   NOR2_X0_50_SVT g45180 (.A(n_22),
	.B(n_16),
	.Q(n_74));
   NAND2_X0_50_SVT g45181 (.A(n_27),
	.B(n_15),
	.Q(n_73));
   NAND2_X4_50_SVT g45182 (.A(n_25),
	.B(n_15),
	.Q(n_72));
   NOR2_X0_50_SVT g45183 (.A(n_28),
	.B(n_14),
	.Q(n_71));
   NOR2_X0_50_SVT g45184 (.A(n_28),
	.B(n_13),
	.Q(n_70));
   NAND2_X0_50_SVT g45185 (.A(n_25),
	.B(n_1),
	.Q(n_69));
   CLKAND2_X6_50_SVT g45186 (.A(n_25),
	.B(n_12),
	.Q(n_68));
   NAND2_X1_50_SVT g45187 (.A(n_21),
	.B(n_12),
	.Q(n_67));
   CLKAND2_X6_50_SVT g45188 (.A(n_23),
	.B(n_12),
	.Q(n_66));
   CLKAND2_X6_50_SVT g45189 (.A(n_25),
	.B(n_18),
	.Q(n_65));
   NAND2_X0_50_SVT g45190 (.A(n_21),
	.B(n_18),
	.Q(n_64));
   CLKAND2_X6_50_SVT g45191 (.A(n_23),
	.B(n_18),
	.Q(n_63));
   CLKNAND2_X4_50_SVT g45193 (.A(n_21),
	.B(n_1),
	.Q(n_62));
   MUX2_X2_50_SVT g45194 (.A(DPATH_n_2913),
	.B(DPATH_n_2881),
	.Q(n_60),
	.S0(n_11));
   MUX2_X2_50_SVT g45195 (.A(DPATH_n_2894),
	.B(DPATH_n_2862),
	.Q(n_59),
	.S0(n_11));
   MUX2_X2_50_SVT g45196 (.A(DPATH_n_2893),
	.B(DPATH_n_2861),
	.Q(n_58),
	.S0(n_11));
   MUX2_X2_50_SVT g45197 (.A(DPATH_n_2902),
	.B(DPATH_n_2870),
	.Q(n_57),
	.S0(n_11));
   MUX2_X2_50_SVT g45198 (.A(DPATH_n_2911),
	.B(DPATH_n_2879),
	.Q(n_56),
	.S0(n_11));
   MUX2_X2_50_SVT g45199 (.A(DPATH_n_2901),
	.B(DPATH_n_2869),
	.Q(n_55),
	.S0(n_11));
   MUX2_X2_50_SVT g45200 (.A(DPATH_n_2899),
	.B(DPATH_n_2867),
	.Q(n_54),
	.S0(n_11));
   MUX2_X2_50_SVT g45202 (.A(DPATH_n_2912),
	.B(DPATH_n_2880),
	.Q(n_52),
	.S0(n_11));
   MUX2_X2_50_SVT g45203 (.A(DPATH_n_2918),
	.B(DPATH_n_2886),
	.Q(n_51),
	.S0(n_11));
   MUX2_X2_50_SVT g45204 (.A(DPATH_n_2917),
	.B(DPATH_n_2885),
	.Q(n_50),
	.S0(n_11));
   MUX2_X2_50_SVT g45205 (.A(DPATH_n_2914),
	.B(DPATH_n_2882),
	.Q(n_49),
	.S0(n_11));
   MUX2_X2_50_SVT g45206 (.A(DPATH_n_2915),
	.B(DPATH_n_2883),
	.Q(n_48),
	.S0(n_11));
   MUX2_X2_50_SVT g45207 (.A(DPATH_n_2907),
	.B(DPATH_n_2875),
	.Q(n_47),
	.S0(n_11));
   MUX2_X2_50_SVT g45208 (.A(DPATH_n_2898),
	.B(DPATH_n_2866),
	.Q(n_46),
	.S0(n_11));
   MUX2_X2_50_SVT g45209 (.A(DPATH_n_2916),
	.B(DPATH_n_2884),
	.Q(n_45),
	.S0(n_11));
   NAND2_A_OAI21_X2_50_SVT g45210 (.A0N(n_10),
	.A1N(DPATH_n_2922),
	.B0(n_10),
	.B1(PC[2]),
	.Q(n_44));
   MUX2_X2_50_SVT g45211 (.A(DPATH_n_2908),
	.B(DPATH_n_2876),
	.Q(n_43),
	.S0(n_11));
   MUX2_X2_50_SVT g45212 (.A(DPATH_n_2920),
	.B(DPATH_n_2888),
	.Q(n_42),
	.S0(n_11));
   MUX2_X2_50_SVT g45213 (.A(DPATH_n_2921),
	.B(DPATH_n_2889),
	.Q(n_41),
	.S0(n_11));
   MUX2_X2_50_SVT g45214 (.A(DPATH_n_2923),
	.B(PC[1]),
	.Q(n_40),
	.S0(n_11));
   MUX2_X2_50_SVT g45215 (.A(DPATH_n_2903),
	.B(DPATH_n_2871),
	.Q(n_39),
	.S0(n_11));
   MUX2_X2_50_SVT g45216 (.A(DPATH_n_2910),
	.B(DPATH_n_2878),
	.Q(n_38),
	.S0(n_11));
   MUX2_X2_50_SVT g45217 (.A(DPATH_n_2895),
	.B(DPATH_n_2863),
	.Q(n_37),
	.S0(n_11));
   MUX2_X2_50_SVT g45218 (.A(DPATH_n_2905),
	.B(DPATH_n_2873),
	.Q(n_36),
	.S0(n_11));
   MUX2_X2_50_SVT g45219 (.A(DPATH_n_2909),
	.B(DPATH_n_2877),
	.Q(n_35),
	.S0(n_11));
   MUX2_X2_50_SVT g45220 (.A(DPATH_n_2897),
	.B(DPATH_n_2865),
	.Q(n_34),
	.S0(n_11));
   MUX2_X2_50_SVT g45221 (.A(DPATH_n_2900),
	.B(DPATH_n_2868),
	.Q(n_33),
	.S0(n_11));
   MUX2_X2_50_SVT g45222 (.A(DPATH_n_2919),
	.B(DPATH_n_2887),
	.Q(n_32),
	.S0(n_11));
   MUX2_X2_50_SVT g45223 (.A(DPATH_n_2904),
	.B(DPATH_n_2872),
	.Q(n_31),
	.S0(n_11));
   MUX2_X2_50_SVT g45224 (.A(DPATH_n_2896),
	.B(DPATH_n_2864),
	.Q(n_30),
	.S0(n_11));
   MUX2_X2_50_SVT g45225 (.A(DPATH_n_2906),
	.B(DPATH_n_2874),
	.Q(n_29),
	.S0(n_11));
   INV_A_NAND2_X0_50_SVT g45228 (.AN(INSTR[8]),
	.B(n_20),
	.Q(n_28));
   NAND2_X0_50_SVT g45229 (.A(n_19),
	.B(INSTR[8]),
	.Q(n_26));
   INV_X2_50_SVT g45231 (.A(n_22),
	.Q(n_21));
   NAND2_X0_50_SVT g45232 (.A(n_20),
	.B(INSTR[8]),
	.Q(n_24));
   INV_A_NAND2_X0_50_SVT g45233 (.AN(INSTR[8]),
	.B(n_19),
	.Q(n_22));
   NOR2_X0_50_SVT g45234 (.A(INSTR[9]),
	.B(n_2835),
	.Q(n_20));
   INV_A_NOR2_X0_50_SVT g45235 (.AN(INSTR[9]),
	.B(n_2835),
	.Q(n_19));
   INV_A_NOR2_X0_50_SVT g45236 (.AN(n_6),
	.B(INSTR[7]),
	.Q(n_18));
   NOR2P3_X1_50_SVT g45237 (.A(INSTR[7]),
	.B(n_9),
	.Q(n_17));
   NAND2T_X0_50_SVT g45238 (.A(n_6),
	.B(INSTR[7]),
	.Q(n_16));
   NOR2P3_X1_50_SVT g45239 (.A(INSTR[7]),
	.B(n_5),
	.Q(n_15));
   INVP2_X1_50_SVT g45241 (.A(n_11),
	.Q(n_10));
   NAND2T_X0_50_SVT g45242 (.A(n_7),
	.B(INSTR[7]),
	.Q(n_14));
   INV_A_NAND2_X0_50_SVT g45243 (.AN(n_5),
	.B(INSTR[7]),
	.Q(n_13));
   INV_A_NOR2_X0_50_SVT g45244 (.AN(INSTR[7]),
	.B(n_9),
	.Q(n_12));
   OA21_X4_50_SVT g45247 (.A0(n_2834),
	.A1(n_2706),
	.B0(n_3),
	.Q(n_11));
   NAND2_X0_50_SVT g45249 (.A(INSTR[10]),
	.B(INSTR[11]),
	.Q(n_9));
   INV_A_NOR2_X0_50_SVT g45251 (.AN(INSTR[10]),
	.B(INSTR[11]),
	.Q(n_7));
   NOR2_X0_50_SVT g45253 (.A(INSTR[10]),
	.B(INSTR[11]),
	.Q(n_6));
   INV_A_NAND2_X0_50_SVT g45254 (.AN(INSTR[10]),
	.B(INSTR[11]),
	.Q(n_5));
   NOR2P3T_X2_50_SVT g45255 (.A(INSTR[5]),
	.B(INSTR[4]),
	.Q(n_4));
   INV_A_NAND2_X0_50_SVT g79925 (.AN(n_28),
	.B(n_12),
	.Q(n_2));
   INV_A_NOR2_X2_50_SVT g45266 (.AN(n_7),
	.B(INSTR[7]),
	.Q(n_1));
   INV_A_NOR2_X4_50_SVT g45267 (.AN(n_3),
	.B(n_4),
	.Q(n_0));
   XOR3_X2_50_SVT DPATH_addinc_ALU_add_381_20_g2274 (.A(DPATH_A_31_),
	.B(n_1149),
	.C(DPATH_addinc_ALU_add_381_20_n_1104),
	.Q(DPATH_ALU_SUM_31__624));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2275 (.A(DPATH_n_2384),
	.B(n_2684),
	.CI(DPATH_addinc_ALU_add_381_20_n_1106),
	.CO(DPATH_addinc_ALU_add_381_20_n_1104),
	.S(DPATH_n_2567));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2276 (.A(DPATH_n_2385),
	.B(n_2677),
	.CI(DPATH_addinc_ALU_add_381_20_n_1108),
	.CO(DPATH_addinc_ALU_add_381_20_n_1106),
	.S(DPATH_n_2568));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2277 (.A(DPATH_n_2386),
	.B(n_2697),
	.CI(DPATH_addinc_ALU_add_381_20_n_1110),
	.CO(DPATH_addinc_ALU_add_381_20_n_1108),
	.S(DPATH_n_2569));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2278 (.A(DPATH_n_2387),
	.B(n_2694),
	.CI(DPATH_addinc_ALU_add_381_20_n_1112),
	.CO(DPATH_addinc_ALU_add_381_20_n_1110),
	.S(DPATH_n_2570));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2279 (.A(DPATH_n_2388),
	.B(n_2683),
	.CI(DPATH_addinc_ALU_add_381_20_n_1114),
	.CO(DPATH_addinc_ALU_add_381_20_n_1112),
	.S(DPATH_n_2571));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2280 (.A(DPATH_n_2389),
	.B(n_2701),
	.CI(DPATH_addinc_ALU_add_381_20_n_1116),
	.CO(DPATH_addinc_ALU_add_381_20_n_1114),
	.S(DPATH_n_2572));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2281 (.A(DPATH_n_2390),
	.B(n_2692),
	.CI(DPATH_addinc_ALU_add_381_20_n_1118),
	.CO(DPATH_addinc_ALU_add_381_20_n_1116),
	.S(DPATH_n_2573));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2282 (.A(DPATH_n_2391),
	.B(n_2703),
	.CI(DPATH_addinc_ALU_add_381_20_n_1120),
	.CO(DPATH_addinc_ALU_add_381_20_n_1118),
	.S(DPATH_n_2574));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2283 (.A(DPATH_n_2392),
	.B(n_2690),
	.CI(DPATH_addinc_ALU_add_381_20_n_1122),
	.CO(DPATH_addinc_ALU_add_381_20_n_1120),
	.S(DPATH_n_2575));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2284 (.A(DPATH_n_2393),
	.B(n_2685),
	.CI(DPATH_addinc_ALU_add_381_20_n_1124),
	.CO(DPATH_addinc_ALU_add_381_20_n_1122),
	.S(DPATH_n_2576));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2285 (.A(DPATH_n_2394),
	.B(n_2682),
	.CI(DPATH_addinc_ALU_add_381_20_n_1126),
	.CO(DPATH_addinc_ALU_add_381_20_n_1124),
	.S(DPATH_n_2577));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2286 (.A(DPATH_n_2395),
	.B(n_2704),
	.CI(DPATH_addinc_ALU_add_381_20_n_1128),
	.CO(DPATH_addinc_ALU_add_381_20_n_1126),
	.S(DPATH_n_2578));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2287 (.A(DPATH_n_2396),
	.B(n_2696),
	.CI(DPATH_addinc_ALU_add_381_20_n_1130),
	.CO(DPATH_addinc_ALU_add_381_20_n_1128),
	.S(DPATH_n_2579));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2288 (.A(DPATH_n_2397),
	.B(n_2695),
	.CI(DPATH_addinc_ALU_add_381_20_n_1132),
	.CO(DPATH_addinc_ALU_add_381_20_n_1130),
	.S(DPATH_n_2580));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2289 (.A(DPATH_n_2398),
	.B(n_2691),
	.CI(DPATH_addinc_ALU_add_381_20_n_1134),
	.CO(DPATH_addinc_ALU_add_381_20_n_1132),
	.S(DPATH_n_2581));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2290 (.A(DPATH_n_2399),
	.B(n_2673),
	.CI(DPATH_addinc_ALU_add_381_20_n_1136),
	.CO(DPATH_addinc_ALU_add_381_20_n_1134),
	.S(DPATH_n_2582));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2291 (.A(DPATH_n_2400),
	.B(n_2686),
	.CI(DPATH_addinc_ALU_add_381_20_n_1138),
	.CO(DPATH_addinc_ALU_add_381_20_n_1136),
	.S(DPATH_n_2583));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2292 (.A(DPATH_n_2401),
	.B(n_2681),
	.CI(DPATH_addinc_ALU_add_381_20_n_1140),
	.CO(DPATH_addinc_ALU_add_381_20_n_1138),
	.S(DPATH_n_2584));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2293 (.A(DPATH_n_2402),
	.B(n_2680),
	.CI(DPATH_addinc_ALU_add_381_20_n_1142),
	.CO(DPATH_addinc_ALU_add_381_20_n_1140),
	.S(DPATH_n_2585));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2294 (.A(DPATH_n_2403),
	.B(n_2678),
	.CI(DPATH_addinc_ALU_add_381_20_n_1144),
	.CO(DPATH_addinc_ALU_add_381_20_n_1142),
	.S(DPATH_n_2586));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2295 (.A(DPATH_n_2404),
	.B(n_2676),
	.CI(DPATH_addinc_ALU_add_381_20_n_1146),
	.CO(DPATH_addinc_ALU_add_381_20_n_1144),
	.S(DPATH_n_2587));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2296 (.A(DPATH_n_2405),
	.B(n_2674),
	.CI(DPATH_addinc_ALU_add_381_20_n_1148),
	.CO(DPATH_addinc_ALU_add_381_20_n_1146),
	.S(DPATH_n_2588));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2297 (.A(DPATH_n_2406),
	.B(n_2688),
	.CI(DPATH_addinc_ALU_add_381_20_n_1150),
	.CO(DPATH_addinc_ALU_add_381_20_n_1148),
	.S(DPATH_n_2589));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2298 (.A(DPATH_n_2407),
	.B(n_2689),
	.CI(DPATH_addinc_ALU_add_381_20_n_1152),
	.CO(DPATH_addinc_ALU_add_381_20_n_1150),
	.S(DPATH_n_2590));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2299 (.A(DPATH_n_2408),
	.B(n_2699),
	.CI(DPATH_addinc_ALU_add_381_20_n_1154),
	.CO(DPATH_addinc_ALU_add_381_20_n_1152),
	.S(DPATH_n_2591));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2300 (.A(DPATH_n_2409),
	.B(n_2679),
	.CI(DPATH_addinc_ALU_add_381_20_n_1156),
	.CO(DPATH_addinc_ALU_add_381_20_n_1154),
	.S(DPATH_n_2592));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2301 (.A(DPATH_n_2410),
	.B(n_2675),
	.CI(DPATH_addinc_ALU_add_381_20_n_1158),
	.CO(DPATH_addinc_ALU_add_381_20_n_1156),
	.S(DPATH_n_2593));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2302 (.A(DPATH_n_2411),
	.B(n_2698),
	.CI(DPATH_addinc_ALU_add_381_20_n_1160),
	.CO(DPATH_addinc_ALU_add_381_20_n_1158),
	.S(DPATH_n_2594));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2303 (.A(DPATH_n_2412),
	.B(n_2693),
	.CI(DPATH_addinc_ALU_add_381_20_n_1162),
	.CO(DPATH_addinc_ALU_add_381_20_n_1160),
	.S(DPATH_n_2595));
   FA1_X1_50_SVT DPATH_addinc_ALU_add_381_20_g2304 (.A(DPATH_n_2413),
	.B(n_2687),
	.CI(DPATH_addinc_ALU_add_381_20_n_1165),
	.CO(DPATH_addinc_ALU_add_381_20_n_1162),
	.S(DPATH_n_2596));
   NAND2_A_NAND2_X2_50_SVT DPATH_addinc_ALU_add_381_20_g2305 (.A0N(n_2702),
	.A1N(DPATH_n_2414),
	.B0(DPATH_addinc_ALU_add_381_20_n_1165),
	.Q(DPATH_n_2597));
   OR2_X2_50_SVT DPATH_addinc_ALU_add_381_20_g2306 (.A(n_2702),
	.B(DPATH_n_2414),
	.Q(DPATH_addinc_ALU_add_381_20_n_1165));
   XOR3_X0_50_SVT DPATH_ADDBRANCH_add_422_17_g750 (.A(PC[31]),
	.B(INSTR[31]),
	.C(DPATH_ADDBRANCH_add_422_17_n_596),
	.Q(DPATH_n_2893));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g751 (.A(INSTR[31]),
	.B(PC[30]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_599),
	.CO(DPATH_ADDBRANCH_add_422_17_n_596),
	.S(DPATH_n_2894));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g752 (.A(INSTR[31]),
	.B(PC[29]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_601),
	.CO(DPATH_ADDBRANCH_add_422_17_n_599),
	.S(DPATH_n_2895));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g753 (.A(INSTR[31]),
	.B(PC[28]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_603),
	.CO(DPATH_ADDBRANCH_add_422_17_n_601),
	.S(DPATH_n_2896));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g754 (.A(INSTR[31]),
	.B(PC[27]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_605),
	.CO(DPATH_ADDBRANCH_add_422_17_n_603),
	.S(DPATH_n_2897));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g755 (.A(INSTR[31]),
	.B(PC[26]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_607),
	.CO(DPATH_ADDBRANCH_add_422_17_n_605),
	.S(DPATH_n_2898));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g756 (.A(INSTR[31]),
	.B(PC[25]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_609),
	.CO(DPATH_ADDBRANCH_add_422_17_n_607),
	.S(DPATH_n_2899));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g757 (.A(INSTR[31]),
	.B(PC[24]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_611),
	.CO(DPATH_ADDBRANCH_add_422_17_n_609),
	.S(DPATH_n_2900));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g758 (.A(INSTR[31]),
	.B(PC[23]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_613),
	.CO(DPATH_ADDBRANCH_add_422_17_n_611),
	.S(DPATH_n_2901));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g759 (.A(INSTR[31]),
	.B(PC[22]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_615),
	.CO(DPATH_ADDBRANCH_add_422_17_n_613),
	.S(DPATH_n_2902));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g760 (.A(INSTR[31]),
	.B(PC[21]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_617),
	.CO(DPATH_ADDBRANCH_add_422_17_n_615),
	.S(DPATH_n_2903));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g761 (.A(INSTR[31]),
	.B(PC[20]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_619),
	.CO(DPATH_ADDBRANCH_add_422_17_n_617),
	.S(DPATH_n_2904));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g762 (.A(DPATH_n_5211),
	.B(PC[19]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_621),
	.CO(DPATH_ADDBRANCH_add_422_17_n_619),
	.S(DPATH_n_2905));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g763 (.A(DPATH_n_5212),
	.B(PC[18]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_623),
	.CO(DPATH_ADDBRANCH_add_422_17_n_621),
	.S(DPATH_n_2906));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g764 (.A(DPATH_n_5213),
	.B(PC[17]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_625),
	.CO(DPATH_ADDBRANCH_add_422_17_n_623),
	.S(DPATH_n_2907));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g765 (.A(DPATH_n_5214),
	.B(PC[16]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_627),
	.CO(DPATH_ADDBRANCH_add_422_17_n_625),
	.S(DPATH_n_2908));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g766 (.A(DPATH_n_5215),
	.B(PC[15]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_629),
	.CO(DPATH_ADDBRANCH_add_422_17_n_627),
	.S(DPATH_n_2909));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g767 (.A(DPATH_n_5216),
	.B(PC[14]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_631),
	.CO(DPATH_ADDBRANCH_add_422_17_n_629),
	.S(DPATH_n_2910));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g768 (.A(DPATH_n_5217),
	.B(PC[13]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_633),
	.CO(DPATH_ADDBRANCH_add_422_17_n_631),
	.S(DPATH_n_2911));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g769 (.A(DPATH_n_5218),
	.B(PC[12]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_635),
	.CO(DPATH_ADDBRANCH_add_422_17_n_633),
	.S(DPATH_n_2912));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g770 (.A(n_2836),
	.B(PC[11]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_637),
	.CO(DPATH_ADDBRANCH_add_422_17_n_635),
	.S(DPATH_n_2913));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g771 (.A(INSTR[30]),
	.B(PC[10]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_639),
	.CO(DPATH_ADDBRANCH_add_422_17_n_637),
	.S(DPATH_n_2914));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g772 (.A(INSTR[29]),
	.B(PC[9]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_641),
	.CO(DPATH_ADDBRANCH_add_422_17_n_639),
	.S(DPATH_n_2915));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g773 (.A(INSTR[28]),
	.B(PC[8]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_643),
	.CO(DPATH_ADDBRANCH_add_422_17_n_641),
	.S(DPATH_n_2916));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g774 (.A(INSTR[27]),
	.B(PC[7]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_645),
	.CO(DPATH_ADDBRANCH_add_422_17_n_643),
	.S(DPATH_n_2917));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g775 (.A(INSTR[26]),
	.B(PC[6]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_647),
	.CO(DPATH_ADDBRANCH_add_422_17_n_645),
	.S(DPATH_n_2918));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g776 (.A(INSTR[25]),
	.B(PC[5]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_649),
	.CO(DPATH_ADDBRANCH_add_422_17_n_647),
	.S(DPATH_n_2919));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g777 (.A(DPATH_n_5226),
	.B(PC[4]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_651),
	.CO(DPATH_ADDBRANCH_add_422_17_n_649),
	.S(DPATH_n_2920));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g778 (.A(DPATH_n_5227),
	.B(PC[3]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_653),
	.CO(DPATH_ADDBRANCH_add_422_17_n_651),
	.S(DPATH_n_2921));
   FA1_X1_50_SVT DPATH_ADDBRANCH_add_422_17_g779 (.A(DPATH_n_5228),
	.B(PC[2]),
	.CI(DPATH_ADDBRANCH_add_422_17_n_655),
	.CO(DPATH_ADDBRANCH_add_422_17_n_653),
	.S(DPATH_n_2922));
   XOR2NG_X1P5_50_SVT DPATH_ADDFOUR_add_172_17_g916 (.A(PC[31]),
	.B(DPATH_ADDFOUR_add_172_17_n_635),
	.Q(DPATH_n_2861));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g917 (.A(PC[30]),
	.B(DPATH_ADDFOUR_add_172_17_n_637),
	.CO(DPATH_ADDFOUR_add_172_17_n_635),
	.S(DPATH_n_2862));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g918 (.A(PC[29]),
	.B(DPATH_ADDFOUR_add_172_17_n_639),
	.CO(DPATH_ADDFOUR_add_172_17_n_637),
	.S(DPATH_n_2863));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g919 (.A(PC[28]),
	.B(DPATH_ADDFOUR_add_172_17_n_641),
	.CO(DPATH_ADDFOUR_add_172_17_n_639),
	.S(DPATH_n_2864));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g920 (.A(PC[27]),
	.B(DPATH_ADDFOUR_add_172_17_n_643),
	.CO(DPATH_ADDFOUR_add_172_17_n_641),
	.S(DPATH_n_2865));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g921 (.A(PC[26]),
	.B(DPATH_ADDFOUR_add_172_17_n_645),
	.CO(DPATH_ADDFOUR_add_172_17_n_643),
	.S(DPATH_n_2866));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g922 (.A(PC[25]),
	.B(DPATH_ADDFOUR_add_172_17_n_647),
	.CO(DPATH_ADDFOUR_add_172_17_n_645),
	.S(DPATH_n_2867));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g923 (.A(PC[24]),
	.B(DPATH_ADDFOUR_add_172_17_n_649),
	.CO(DPATH_ADDFOUR_add_172_17_n_647),
	.S(DPATH_n_2868));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g924 (.A(PC[23]),
	.B(DPATH_ADDFOUR_add_172_17_n_651),
	.CO(DPATH_ADDFOUR_add_172_17_n_649),
	.S(DPATH_n_2869));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g925 (.A(PC[22]),
	.B(DPATH_ADDFOUR_add_172_17_n_653),
	.CO(DPATH_ADDFOUR_add_172_17_n_651),
	.S(DPATH_n_2870));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g926 (.A(PC[21]),
	.B(DPATH_ADDFOUR_add_172_17_n_655),
	.CO(DPATH_ADDFOUR_add_172_17_n_653),
	.S(DPATH_n_2871));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g927 (.A(PC[20]),
	.B(DPATH_ADDFOUR_add_172_17_n_657),
	.CO(DPATH_ADDFOUR_add_172_17_n_655),
	.S(DPATH_n_2872));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g928 (.A(PC[19]),
	.B(DPATH_ADDFOUR_add_172_17_n_659),
	.CO(DPATH_ADDFOUR_add_172_17_n_657),
	.S(DPATH_n_2873));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g929 (.A(PC[18]),
	.B(DPATH_ADDFOUR_add_172_17_n_661),
	.CO(DPATH_ADDFOUR_add_172_17_n_659),
	.S(DPATH_n_2874));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g930 (.A(PC[17]),
	.B(DPATH_ADDFOUR_add_172_17_n_663),
	.CO(DPATH_ADDFOUR_add_172_17_n_661),
	.S(DPATH_n_2875));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g931 (.A(PC[16]),
	.B(DPATH_ADDFOUR_add_172_17_n_665),
	.CO(DPATH_ADDFOUR_add_172_17_n_663),
	.S(DPATH_n_2876));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g932 (.A(PC[15]),
	.B(DPATH_ADDFOUR_add_172_17_n_667),
	.CO(DPATH_ADDFOUR_add_172_17_n_665),
	.S(DPATH_n_2877));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g933 (.A(PC[14]),
	.B(DPATH_ADDFOUR_add_172_17_n_669),
	.CO(DPATH_ADDFOUR_add_172_17_n_667),
	.S(DPATH_n_2878));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g934 (.A(PC[13]),
	.B(DPATH_ADDFOUR_add_172_17_n_671),
	.CO(DPATH_ADDFOUR_add_172_17_n_669),
	.S(DPATH_n_2879));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g935 (.A(PC[12]),
	.B(DPATH_ADDFOUR_add_172_17_n_673),
	.CO(DPATH_ADDFOUR_add_172_17_n_671),
	.S(DPATH_n_2880));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g936 (.A(PC[11]),
	.B(DPATH_ADDFOUR_add_172_17_n_675),
	.CO(DPATH_ADDFOUR_add_172_17_n_673),
	.S(DPATH_n_2881));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g937 (.A(PC[10]),
	.B(DPATH_ADDFOUR_add_172_17_n_677),
	.CO(DPATH_ADDFOUR_add_172_17_n_675),
	.S(DPATH_n_2882));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g938 (.A(PC[9]),
	.B(DPATH_ADDFOUR_add_172_17_n_679),
	.CO(DPATH_ADDFOUR_add_172_17_n_677),
	.S(DPATH_n_2883));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g939 (.A(PC[8]),
	.B(DPATH_ADDFOUR_add_172_17_n_681),
	.CO(DPATH_ADDFOUR_add_172_17_n_679),
	.S(DPATH_n_2884));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g940 (.A(PC[7]),
	.B(DPATH_ADDFOUR_add_172_17_n_683),
	.CO(DPATH_ADDFOUR_add_172_17_n_681),
	.S(DPATH_n_2885));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g941 (.A(PC[6]),
	.B(DPATH_ADDFOUR_add_172_17_n_685),
	.CO(DPATH_ADDFOUR_add_172_17_n_683),
	.S(DPATH_n_2886));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g942 (.A(PC[5]),
	.B(DPATH_ADDFOUR_add_172_17_n_687),
	.CO(DPATH_ADDFOUR_add_172_17_n_685),
	.S(DPATH_n_2887));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g943 (.A(PC[4]),
	.B(DPATH_ADDFOUR_add_172_17_n_689),
	.CO(DPATH_ADDFOUR_add_172_17_n_687),
	.S(DPATH_n_2888));
   HA1_X1_50_SVT DPATH_ADDFOUR_add_172_17_g944 (.A(PC[2]),
	.B(PC[3]),
	.CO(DPATH_ADDFOUR_add_172_17_n_689),
	.S(DPATH_n_2889));
   NAND4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g815 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_58),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_66),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_67),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_70),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_71));
   NOR4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g816 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_55),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_65),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_69),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_63),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_70));
   NAND4T_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g817 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_62),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_40),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_45),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_60),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_69));
   NAND4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g818 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_22),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_43),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_39),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_51),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_68));
   NOR4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g819 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_44),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_53),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_42),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_56),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_67));
   NOR4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g820 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_36),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_34),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_48),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_32),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_66));
   NAND4T_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g821 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_52),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_31),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_35),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_54),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_65));
   NAND4_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g822 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_33),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_49),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_59),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_57),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_64));
   NAND4T_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g823 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_37),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_47),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_61),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_50),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_63));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g824 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_10),
	.B(DPATH_n_2818),
	.C(DPATH_n_2780),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_62));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g825 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_18),
	.B(DPATH_n_2822),
	.C(DPATH_n_2784),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_61));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g826 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_21),
	.B(DPATH_n_2825),
	.C(DPATH_n_2787),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_60));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g827 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_19),
	.B(DPATH_n_2803),
	.C(DPATH_n_2765),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_59));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g828 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_16),
	.B(DPATH_n_2800),
	.C(DPATH_n_2762),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_58));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g829 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_17),
	.B(DPATH_n_2807),
	.C(DPATH_n_2769),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_57));
   XNOR3_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g830 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_9),
	.B(DPATH_n_2814),
	.C(DPATH_n_2776),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_56));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g831 (.A(DPATH_n_2811),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_20),
	.C(DPATH_n_2773),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_55));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g832 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_25),
	.B(DPATH_n_2817),
	.C(DPATH_n_2779),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_54));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g833 (.A(DPATH_n_2810),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_27),
	.C(DPATH_n_2772),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_53));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g834 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_26),
	.B(DPATH_n_2813),
	.C(DPATH_n_2775),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_52));
   XOR3_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g835 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_29),
	.B(DPATH_n_2799),
	.C(DPATH_n_2761),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_51));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g836 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_30),
	.B(DPATH_n_2824),
	.C(DPATH_n_2786),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_50));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g837 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_28),
	.B(DPATH_n_2802),
	.C(DPATH_n_2764),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_49));
   XNOR3_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g838 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_23),
	.B(DPATH_n_2806),
	.C(DPATH_n_2768),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_48));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g839 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_24),
	.B(DPATH_n_2821),
	.C(DPATH_n_2783),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_47));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g840 (.A(DPATH_n_2796),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_4),
	.C(DPATH_n_2758),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_46));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g841 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_38),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_41),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_45));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g842 (.A(DPATH_n_2809),
	.B(DPATH_n_2771),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_0),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_44));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g843 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_7),
	.B(DPATH_n_2797),
	.C(DPATH_n_2759),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_43));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g844 (.A(DPATH_n_2812),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_15),
	.C(DPATH_n_2774),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_42));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g845 (.A(DPATH_n_2823),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_13),
	.C(DPATH_n_2785),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_41));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g846 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_3),
	.B(DPATH_n_2819),
	.C(DPATH_n_2781),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_40));
   XOR3_X1_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g847 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_5),
	.B(DPATH_n_2798),
	.C(DPATH_n_2760),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_39));
   XOR3_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g848 (.A(DPATH_n_2826),
	.B(DPATH_n_2827),
	.C(DPATH_n_2788),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_38));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g849 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_2),
	.B(DPATH_n_2820),
	.C(DPATH_n_2782),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_37));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g850 (.A(DPATH_n_2804),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_8),
	.C(DPATH_n_2766),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_36));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g851 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_14),
	.B(DPATH_n_2816),
	.C(DPATH_n_2778),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_35));
   XNOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g852 (.A(DPATH_n_2805),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_11),
	.C(DPATH_n_2767),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_34));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g853 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_1),
	.B(DPATH_n_2801),
	.C(DPATH_n_2763),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_33));
   XNOR3_X0_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g854 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_12),
	.B(DPATH_n_2808),
	.C(DPATH_n_2770),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_32));
   XOR3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g855 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_6),
	.B(DPATH_n_2815),
	.C(DPATH_n_2777),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_31));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g856 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_21),
	.B(DPATH_n_2825),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_30));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g857 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_16),
	.B(DPATH_n_2800),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_29));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g858 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_19),
	.B(DPATH_n_2803),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_28));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g859 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_20),
	.B(DPATH_n_2811),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_27));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g860 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_9),
	.B(DPATH_n_2814),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_26));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g861 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_10),
	.B(DPATH_n_2818),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_25));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g862 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_18),
	.B(DPATH_n_2822),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_24));
   INV_A_NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g863 (.AN(DPATH_csa_tree_ALU_eq_397_21_groupi_n_17),
	.B(DPATH_n_2807),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_23));
   XNOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g864 (.A(DPATH_n_2789),
	.B(DPATH_n_2827),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_22));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g865 (.A(DPATH_n_2775),
	.B(DPATH_n_2813),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_15));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g866 (.A(DPATH_n_2817),
	.B(DPATH_n_2779),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_14));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g867 (.A(DPATH_n_2824),
	.B(DPATH_n_2786),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_13));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g868 (.A(DPATH_n_2809),
	.B(DPATH_n_2771),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_12));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g869 (.A(DPATH_n_2768),
	.B(DPATH_n_2806),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_11));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g870 (.A(DPATH_n_2827),
	.B(DPATH_n_2826),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_21));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g871 (.A(DPATH_n_2812),
	.B(DPATH_n_2774),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_20));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g872 (.A(DPATH_n_2804),
	.B(DPATH_n_2766),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_19));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g873 (.A(DPATH_n_2823),
	.B(DPATH_n_2785),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_18));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g874 (.A(DPATH_n_2808),
	.B(DPATH_n_2770),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_17));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g875 (.A(DPATH_n_2801),
	.B(DPATH_n_2763),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_16));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g876 (.A(DPATH_n_2767),
	.B(DPATH_n_2805),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_8));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g877 (.A(DPATH_n_2760),
	.B(DPATH_n_2798),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_7));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g878 (.A(DPATH_n_2816),
	.B(DPATH_n_2778),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_6));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g879 (.A(DPATH_n_2761),
	.B(DPATH_n_2799),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_5));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g880 (.A(DPATH_n_2797),
	.B(DPATH_n_2759),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_4));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g881 (.A(DPATH_n_2820),
	.B(DPATH_n_2782),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_3));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g882 (.A(DPATH_n_2821),
	.B(DPATH_n_2783),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_2));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g883 (.A(DPATH_n_2764),
	.B(DPATH_n_2802),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_1));
   NOR2_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g884 (.A(DPATH_n_2772),
	.B(DPATH_n_2810),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_0));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g885 (.A(DPATH_n_2819),
	.B(DPATH_n_2781),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_10));
   NOR2P3_X2_50_SVT DPATH_csa_tree_ALU_eq_397_21_groupi_g886 (.A(DPATH_n_2815),
	.B(DPATH_n_2777),
	.Q(DPATH_csa_tree_ALU_eq_397_21_groupi_n_9));
   HA1_X1_50_SVT g79927 (.A(DPATH_n_5229),
	.B(PC[1]),
	.CO(DPATH_ADDBRANCH_add_422_17_n_655),
	.S(DPATH_n_2923));
   MUX2_X2_50_SVT g79928 (.A(INSTR[20]),
	.B(INSTR[7]),
	.Q(n_2831),
	.S0(n_1468));
   OR4_X2_50_SVT g79931 (.A(DPATH_csa_tree_ALU_eq_397_21_groupi_n_68),
	.B(DPATH_csa_tree_ALU_eq_397_21_groupi_n_46),
	.C(DPATH_csa_tree_ALU_eq_397_21_groupi_n_71),
	.D(DPATH_csa_tree_ALU_eq_397_21_groupi_n_64),
	.Q(n_2834));
   INV_A_NAND2_X2_50_SVT g79932 (.AN(MEMWRITE),
	.B(n_2706),
	.Q(n_2835));
   AO22_X0_50_SVT g79933 (.A0(INSTR[7]),
	.A1(n_1451),
	.B0(INSTR[20]),
	.B1(INSTR[2]),
	.Q(n_2836));
endmodule

