`timescale 1ns/1ps
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Project: RV32I
//Block: MUX3to1
//HDL: SystemVerilog
//Author : Shamil Niftaliyev
//Reference: "Digital Design and Computer Architecture" D.M.Harris & S.L.Harris (Second Edition)
//Revision history:
//V1: September 15, 2024: 
//Short Summary:
// Three to one digital muliplexer
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////// MODULE DECLARATION
module MUX3to1 (A, B, C, S, Q);
// IOs
  input  logic [31:0] A;        // First argument
  input  logic [31:0] B;        // Second argument
  input  logic [31:0] C;        // Third argument
  input  logic [1:0]  S;        // Select signal
  output logic [31:0] Q;        // Result of multiplexing
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////// 
////// ARCHITECTURE
// Main combinational logic    
  always_comb
  case (S)
    2'b00: Q = A;
    2'b01: Q = B;
    2'b10: Q = C;
    2'b11: Q = 32'bx;
  endcase
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////// 
// END 
endmodule
