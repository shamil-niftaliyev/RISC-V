//systemVerilog HDL for "MAD_RISC_tb", "ADD4_tb" "systemVerilog"


module ADD4_tb ( );

endmodule
