//systemVerilog HDL for "MAD_RISC_tb", "PCREG_tb" "systemVerilog"


module PCREG_tb ( );

endmodule
